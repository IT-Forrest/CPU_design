
module SHARE_SUPERALU_VG ( CLK, RST_N, X_IN, Y_IN, ALU_START, ALU_TYPE, MODE_TYPE, 
        OFFSET, FOUT, POUT, ALU_IS_DONE );
  input [12:0] X_IN;
  input [12:0] Y_IN;
  input [2:0] ALU_TYPE;
  input [1:0] MODE_TYPE;
  input [9:0] OFFSET;
  output [12:0] FOUT;
  output [12:0] POUT;
  input CLK, RST_N, ALU_START;
  output ALU_IS_DONE;
  wire   POST_WORK, PRE_WORK, \INDEX[2] , \RSHT_BITS[3] , SIGN_Y, C152_DATA4_0,
         C152_DATA4_1, C152_DATA4_2, C152_DATA4_3, C152_DATA4_4, C152_DATA4_5,
         C152_DATA4_6, C152_DATA4_7, C152_DATA4_8, C152_DATA4_9, C152_DATA4_10,
         C152_DATA4_11, N74, N90, N91, N92, N121, N122, N123, N124, N128, N129,
         N657, N658, N659, N660, N661, N662, N663, N664, N665, N666, N667,
         N668, N669, N670, N671, N672, N673, N674, N675, N676, N677, N678,
         N679, N680, N681, N682, N683, N684, N685, N686, N687, N688, N689,
         N690, N691, N692, N693, N694, N695, N696, N697, N698, N699, N700,
         N701, N702, N703, N704, N705, N706, N707, N708, N709, N710, N711,
         N712, N713, N714, N715, N716, N717, N718, N719, N720, N721, N722,
         N723, N724, N725, N726, C2_Z_11, C2_Z_10, C2_Z_9, C2_Z_8, C2_Z_7,
         C2_Z_6, C2_Z_5, C2_Z_4, C2_Z_3, C2_Z_2, C2_Z_1, C2_Z_0,
         DP_OP_333_124_4748_N57, DP_OP_333_124_4748_N29,
         DP_OP_333_124_4748_N28, DP_OP_333_124_4748_N27,
         DP_OP_333_124_4748_N26, DP_OP_333_124_4748_N25,
         DP_OP_333_124_4748_N24, DP_OP_333_124_4748_N23,
         DP_OP_333_124_4748_N22, DP_OP_333_124_4748_N21,
         DP_OP_333_124_4748_N20, DP_OP_333_124_4748_N19,
         DP_OP_333_124_4748_N18, DP_OP_333_124_4748_N12,
         DP_OP_333_124_4748_N11, DP_OP_333_124_4748_N10, DP_OP_333_124_4748_N9,
         DP_OP_333_124_4748_N8, DP_OP_333_124_4748_N7, DP_OP_333_124_4748_N6,
         DP_OP_333_124_4748_N5, DP_OP_333_124_4748_N4, DP_OP_333_124_4748_N3,
         DP_OP_333_124_4748_N2, DP_OP_333_124_4748_N1, INTADD_0_CI,
         \INTADD_0_SUM[6] , \INTADD_0_SUM[5] , \INTADD_0_SUM[4] ,
         \INTADD_0_SUM[3] , \INTADD_0_SUM[2] , \INTADD_0_SUM[1] ,
         \INTADD_0_SUM[0] , INTADD_0_N7, INTADD_0_N6, INTADD_0_N5, INTADD_0_N4,
         INTADD_0_N3, INTADD_0_N2, INTADD_0_N1, ADD_X_132_1_N13,
         ADD_X_132_1_N12, ADD_X_132_1_N11, ADD_X_132_1_N10, ADD_X_132_1_N9,
         ADD_X_132_1_N8, ADD_X_132_1_N7, ADD_X_132_1_N6, ADD_X_132_1_N5,
         ADD_X_132_1_N4, ADD_X_132_1_N3, ADD_X_132_1_N2, N1, N2, N3, N4, N5,
         N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N65, N84, N85, N86, N87, N88, N89, N93, N94, N95, N96, N97, N98,
         N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N125,
         N126, N127, N130, N131, N132, N133, N134, N135, N136, N137, N138,
         N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149,
         N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160,
         N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171,
         N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182,
         N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193,
         N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204,
         N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215,
         N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226,
         N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237,
         N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248,
         N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259,
         N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270,
         N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281,
         N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292,
         N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303,
         N304, N305, N306, N307, N308, N309, N310, N311, N312, N313, N314,
         N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325,
         N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336,
         N337, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347,
         N348, N349, N350, N351, N352, N353, N354, N355, N356, N357, N358,
         N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, N369,
         N370, N371, N372, N373, N374, N375, N376, N377, N378, N379, N380,
         N381, N382, N383, N384, N385, N386, N387, N388, N389, N390, N391,
         N392, N393, N394, N395, N396, N397, N398, N399, N400, N401, N402,
         N403, N404, N405, N406, N407, N408, N409, N410, N411, N412, N413,
         N414, N415, N416, N417, N418, N419, N420, N421, N422, N423, N424,
         N425, N426, N427, N428, N429, N430, N431, N432, N433, N434, N435,
         N436, N437, N438, N439, N440, N441, N442, N443, N444, N445, N446,
         N447, N448, N449, N450, N451, N452, N453, N454, N455, N456, N457,
         N458, N459, N460, N461, N462, N463, N464, N465, N466, N467, N468,
         N469, N470, N471, N472, N473, N474, N475, N476, N477, N478, N479,
         N480, N481, N482, N483, N484, N485, N486, N487, N488, N489, N490,
         N491, N492, N493, N494, N495, N496, N497, N498, N499, N500, N501,
         N502, N503, N504, N505, N506, N507, N508, N509, N510, N511, N512,
         N513, N514, N515, N516, N517, N518, N519, N520, N521, N522, N523,
         N524, N525, N526, N527, N528, N529, N530, N531, N532, N533, N534,
         N535, N536, N537, N538, N539, N540, N541, N542, N543, N544, N545,
         N546, N547, N548, N549, N550, N551, N552, N553, N554, N555, N556,
         N557, N558, N559, N560, N561, N562, N563, N564, N565, N566, N567,
         N568, N569, N570, N571, N572, N573, N574, N575, N576, N577, N578,
         N579, N580, N581, N582, N583, N584, N585, N586, N587, N588, N589,
         N590, N591, N592, N593, N594, N595, N596, N597, N598, N599, N600,
         N601, N602, N603, N604, N605, N606, N607, N608, N609, N610, N611,
         N612, N613, N614, N615, N616, N617, N618, N619, N620, N621, N622,
         N623, N624, N625, N626, N627, N628, N629, N630, N631, N632, N633,
         N634, N635, N636, N637, N638, N639, N640, N641, N642, N643, N644,
         N645, N646, N647, N648, N649, N650, N651, N652, N653, N654, N655,
         N656, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736,
         N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747,
         N748, N749, N750, N751, N752, N753, N754, N755, N756, N757, N758,
         N759, N760, N761, N762, N763, N764, N765, N766, N767, N768, N769,
         N770, N771, N772, N773, N774, N775, N776, N777, N778, N779, N780,
         N781, N782, N783, N784, N785, N786, N787, N788, N789, N790, N791,
         N792, N793, N794, N795, N796, N797, N798, N799, N800, N801, N802,
         N803, N804, N805, N806, N807, N808, N809, N810, N811, N812, N813,
         N814, N815, N816, N817, N818, N819, N820, N821, N822, N823, N824,
         N825, N826, N827, N828, N829, N830, N831, N832, N833, N834, N835,
         N836, N837, N838, N839, N840, N841, N842, N843, N844, N845, N846,
         N847, N848, N849, N850, N851, N852, N853, N854, N855, N856, N857,
         N858, N859, N860, N861, N862, N863, N864, N865, N866, N867, N868,
         N869, N870, N871, N872, N873, N874, N875, N876, N877, N878, N879,
         N880, N881, N882, N883, N884, N885, N886, N887, N888, N889, N890,
         N891, N892, N893, N894, N895, N896, N897, N898, N899, N900, N901,
         N902, N903, N904, N905, N906, N907, N908, N909, N910, N911, N912,
         N913, N914, N915, N916, N917, N918, N919, N920, N921, N922, N923,
         N924, N925, N926, N927, N928, N929, N930, N931, N932, N933, N934,
         N935, N936, N937, N938, N939, N940, N941, N942, N943, N944, N945,
         N946, N947, N948, N949, N950, N951, N952, N953, N954, N955, N956,
         N957, N958, N959, N960, N961, N962, N963, N964, N965, N966, N967,
         N968, N969, N970, N971, N972, N973, N974, N975, N976, N977, N978,
         N979, N980, N981, N982, N983, N984, N985, N986, N987, N988, N989,
         N990, N991, N992, N993, N994, N995, N996, N997, N998, N999, N1000,
         N1001, N1002, N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010,
         N1011, N1012, N1013, N1014, N1015;
  wire   [12:9] XTEMP;
  wire   [12:0] DIVISION_HEAD;
  wire   [8:0] DIVISION_REMA;
  wire   [12:0] OPER_A;
  wire   [12:0] OPER_B;
  wire   [12:0] SUM_AB;
  wire   [12:0] ZTEMP;
  wire   [3:2] STEP;

  XOR2X1TF \DP_OP_333_124_4748/U28  ( .A(N85), .B(C2_Z_0), .Y(
        DP_OP_333_124_4748_N29) );
  XOR2X1TF \DP_OP_333_124_4748/U27  ( .A(N85), .B(C2_Z_1), .Y(
        DP_OP_333_124_4748_N28) );
  XOR2X1TF \DP_OP_333_124_4748/U26  ( .A(N85), .B(C2_Z_2), .Y(
        DP_OP_333_124_4748_N27) );
  XOR2X1TF \DP_OP_333_124_4748/U25  ( .A(N85), .B(C2_Z_3), .Y(
        DP_OP_333_124_4748_N26) );
  XOR2X1TF \DP_OP_333_124_4748/U24  ( .A(N967), .B(C2_Z_4), .Y(
        DP_OP_333_124_4748_N25) );
  XOR2X1TF \DP_OP_333_124_4748/U23  ( .A(N85), .B(C2_Z_5), .Y(
        DP_OP_333_124_4748_N24) );
  XOR2X1TF \DP_OP_333_124_4748/U22  ( .A(N967), .B(C2_Z_6), .Y(
        DP_OP_333_124_4748_N23) );
  XOR2X1TF \DP_OP_333_124_4748/U21  ( .A(N85), .B(C2_Z_7), .Y(
        DP_OP_333_124_4748_N22) );
  XOR2X1TF \DP_OP_333_124_4748/U20  ( .A(N967), .B(C2_Z_8), .Y(
        DP_OP_333_124_4748_N21) );
  XOR2X1TF \DP_OP_333_124_4748/U19  ( .A(N85), .B(C2_Z_9), .Y(
        DP_OP_333_124_4748_N20) );
  XOR2X1TF \DP_OP_333_124_4748/U18  ( .A(N967), .B(C2_Z_10), .Y(
        DP_OP_333_124_4748_N19) );
  XOR2X1TF \DP_OP_333_124_4748/U17  ( .A(N85), .B(C2_Z_11), .Y(
        DP_OP_333_124_4748_N18) );
  CMPR32X2TF \DP_OP_333_124_4748/U13  ( .A(DP_OP_333_124_4748_N57), .B(N85), 
        .C(DP_OP_333_124_4748_N29), .CO(DP_OP_333_124_4748_N12), .S(
        C152_DATA4_0) );
  ADDHXLTF \DP_OP_333_124_4748/U12  ( .A(DP_OP_333_124_4748_N28), .B(
        DP_OP_333_124_4748_N12), .CO(DP_OP_333_124_4748_N11), .S(C152_DATA4_1)
         );
  ADDHXLTF \DP_OP_333_124_4748/U11  ( .A(DP_OP_333_124_4748_N27), .B(
        DP_OP_333_124_4748_N11), .CO(DP_OP_333_124_4748_N10), .S(C152_DATA4_2)
         );
  ADDHXLTF \DP_OP_333_124_4748/U10  ( .A(DP_OP_333_124_4748_N26), .B(
        DP_OP_333_124_4748_N10), .CO(DP_OP_333_124_4748_N9), .S(C152_DATA4_3)
         );
  ADDHXLTF \DP_OP_333_124_4748/U9  ( .A(DP_OP_333_124_4748_N25), .B(
        DP_OP_333_124_4748_N9), .CO(DP_OP_333_124_4748_N8), .S(C152_DATA4_4)
         );
  ADDHXLTF \DP_OP_333_124_4748/U8  ( .A(DP_OP_333_124_4748_N24), .B(
        DP_OP_333_124_4748_N8), .CO(DP_OP_333_124_4748_N7), .S(C152_DATA4_5)
         );
  ADDHXLTF \DP_OP_333_124_4748/U7  ( .A(DP_OP_333_124_4748_N23), .B(
        DP_OP_333_124_4748_N7), .CO(DP_OP_333_124_4748_N6), .S(C152_DATA4_6)
         );
  ADDHXLTF \DP_OP_333_124_4748/U6  ( .A(DP_OP_333_124_4748_N22), .B(
        DP_OP_333_124_4748_N6), .CO(DP_OP_333_124_4748_N5), .S(C152_DATA4_7)
         );
  ADDHXLTF \DP_OP_333_124_4748/U5  ( .A(DP_OP_333_124_4748_N21), .B(
        DP_OP_333_124_4748_N5), .CO(DP_OP_333_124_4748_N4), .S(C152_DATA4_8)
         );
  ADDHXLTF \DP_OP_333_124_4748/U4  ( .A(DP_OP_333_124_4748_N20), .B(
        DP_OP_333_124_4748_N4), .CO(DP_OP_333_124_4748_N3), .S(C152_DATA4_9)
         );
  ADDHXLTF \DP_OP_333_124_4748/U3  ( .A(DP_OP_333_124_4748_N19), .B(
        DP_OP_333_124_4748_N3), .CO(DP_OP_333_124_4748_N2), .S(C152_DATA4_10)
         );
  ADDHXLTF \DP_OP_333_124_4748/U2  ( .A(DP_OP_333_124_4748_N18), .B(
        DP_OP_333_124_4748_N2), .CO(DP_OP_333_124_4748_N1), .S(C152_DATA4_11)
         );
  CMPR32X2TF \intadd_0/U8  ( .A(X_IN[1]), .B(DIVISION_HEAD[5]), .C(INTADD_0_CI), .CO(INTADD_0_N7), .S(\INTADD_0_SUM[0] ) );
  CMPR32X2TF \intadd_0/U7  ( .A(X_IN[2]), .B(DIVISION_HEAD[6]), .C(INTADD_0_N7), .CO(INTADD_0_N6), .S(\INTADD_0_SUM[1] ) );
  CMPR32X2TF \intadd_0/U6  ( .A(X_IN[3]), .B(DIVISION_HEAD[7]), .C(INTADD_0_N6), .CO(INTADD_0_N5), .S(\INTADD_0_SUM[2] ) );
  CMPR32X2TF \intadd_0/U5  ( .A(X_IN[4]), .B(DIVISION_HEAD[8]), .C(INTADD_0_N5), .CO(INTADD_0_N4), .S(\INTADD_0_SUM[3] ) );
  CMPR32X2TF \intadd_0/U4  ( .A(X_IN[5]), .B(DIVISION_HEAD[9]), .C(INTADD_0_N4), .CO(INTADD_0_N3), .S(\INTADD_0_SUM[4] ) );
  CMPR32X2TF \intadd_0/U3  ( .A(X_IN[6]), .B(DIVISION_HEAD[10]), .C(
        INTADD_0_N3), .CO(INTADD_0_N2), .S(\INTADD_0_SUM[5] ) );
  CMPR32X2TF \intadd_0/U2  ( .A(X_IN[7]), .B(DIVISION_HEAD[11]), .C(
        INTADD_0_N2), .CO(INTADD_0_N1), .S(\INTADD_0_SUM[6] ) );
  DFFRX2TF \wtemp_reg[3]  ( .D(N679), .CK(CLK), .RN(RST_N), .Q(OPER_B[3]), 
        .QN(N181) );
  DFFSX2TF pre_work_reg ( .D(N695), .CK(CLK), .SN(RST_N), .Q(PRE_WORK), .QN(
        N174) );
  DFFRX2TF \xtemp_reg[10]  ( .D(N709), .CK(CLK), .RN(RST_N), .Q(XTEMP[10]), 
        .QN(N160) );
  DFFRX2TF \ytemp_reg[9]  ( .D(N685), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[0]), .QN(N156) );
  DFFRX2TF \xtemp_reg[11]  ( .D(N708), .CK(CLK), .RN(RST_N), .Q(XTEMP[11]), 
        .QN(N153) );
  DFFRX2TF \xtemp_reg[3]  ( .D(N716), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[7]), .QN(N152) );
  DFFRX2TF \ytemp_reg[10]  ( .D(N684), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[1]), .QN(N149) );
  ADDHX1TF \add_x_132_1/U14  ( .A(OPER_B[0]), .B(OPER_A[0]), .CO(
        ADD_X_132_1_N13), .S(SUM_AB[0]) );
  CMPR32X2TF \add_x_132_1/U4  ( .A(OPER_A[10]), .B(OPER_B[10]), .C(
        ADD_X_132_1_N4), .CO(ADD_X_132_1_N3), .S(SUM_AB[10]) );
  CMPR32X2TF \add_x_132_1/U6  ( .A(OPER_A[8]), .B(OPER_B[8]), .C(
        ADD_X_132_1_N6), .CO(ADD_X_132_1_N5), .S(SUM_AB[8]) );
  CMPR32X2TF \add_x_132_1/U10  ( .A(OPER_A[4]), .B(OPER_B[4]), .C(
        ADD_X_132_1_N10), .CO(ADD_X_132_1_N9), .S(SUM_AB[4]) );
  CMPR32X2TF \add_x_132_1/U12  ( .A(OPER_A[2]), .B(OPER_B[2]), .C(
        ADD_X_132_1_N12), .CO(ADD_X_132_1_N11), .S(SUM_AB[2]) );
  CMPR32X2TF \add_x_132_1/U13  ( .A(OPER_A[1]), .B(OPER_B[1]), .C(
        ADD_X_132_1_N13), .CO(ADD_X_132_1_N12), .S(SUM_AB[1]) );
  CMPR32X2TF \add_x_132_1/U5  ( .A(OPER_A[9]), .B(OPER_B[9]), .C(
        ADD_X_132_1_N5), .CO(ADD_X_132_1_N4), .S(SUM_AB[9]) );
  CMPR32X2TF \add_x_132_1/U11  ( .A(OPER_A[3]), .B(OPER_B[3]), .C(
        ADD_X_132_1_N11), .CO(ADD_X_132_1_N10), .S(SUM_AB[3]) );
  CMPR32X2TF \add_x_132_1/U9  ( .A(OPER_A[5]), .B(OPER_B[5]), .C(
        ADD_X_132_1_N9), .CO(ADD_X_132_1_N8), .S(SUM_AB[5]) );
  CMPR32X2TF \add_x_132_1/U3  ( .A(OPER_A[11]), .B(OPER_B[11]), .C(
        ADD_X_132_1_N3), .CO(ADD_X_132_1_N2), .S(SUM_AB[11]) );
  DFFRX1TF \rsht_bits_reg[2]  ( .D(N701), .CK(CLK), .RN(RST_N), .QN(N90) );
  DFFRX2TF sign_y_reg ( .D(N694), .CK(CLK), .RN(RST_N), .Q(SIGN_Y), .QN(N176)
         );
  DFFRX2TF XOR_SRC_reg ( .D(N707), .CK(CLK), .RN(RST_N), .Q(N63), .QN(N108) );
  DFFRX2TF \rsht_bits_reg[0]  ( .D(N703), .CK(CLK), .RN(RST_N), .Q(N178), .QN(
        N92) );
  DFFRX2TF \step_reg[1]  ( .D(N700), .CK(CLK), .RN(RST_N), .Q(N161), .QN(N121)
         );
  DFFRX2TF \step_reg[3]  ( .D(N721), .CK(CLK), .RN(RST_N), .Q(STEP[3]), .QN(
        N162) );
  DFFRX2TF \step_reg[2]  ( .D(N696), .CK(CLK), .RN(RST_N), .Q(STEP[2]), .QN(
        N150) );
  DFFRX2TF \rsht_bits_reg[1]  ( .D(N702), .CK(CLK), .RN(RST_N), .Q(N167), .QN(
        N91) );
  DFFRX2TF \step_reg[0]  ( .D(N697), .CK(CLK), .RN(RST_N), .Q(N172), .QN(N122)
         );
  DFFRX2TF \rsht_bits_reg[3]  ( .D(N704), .CK(CLK), .RN(RST_N), .Q(
        \RSHT_BITS[3] ), .QN(N187) );
  DFFRX2TF SEL_SRC_reg ( .D(N720), .CK(CLK), .RN(RST_N), .Q(POST_WORK), .QN(
        N171) );
  DFFRX2TF \index_reg[1]  ( .D(N699), .CK(CLK), .RN(RST_N), .Q(N179), .QN(N128) );
  DFFRX2TF SEL_Z_reg ( .D(N670), .CK(CLK), .RN(RST_N), .Q(N173), .QN(N123) );
  DFFRX2TF \index_reg[3]  ( .D(N725), .CK(CLK), .RN(RST_N), .Q(N184), .QN(N124) );
  DFFRX2TF \index_reg[0]  ( .D(N726), .CK(CLK), .RN(RST_N), .Q(N166), .QN(N129) );
  DFFRX2TF \ytemp_reg[0]  ( .D(N705), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[0]), .QN(N177) );
  DFFRX2TF \wtemp_reg[8]  ( .D(N674), .CK(CLK), .RN(RST_N), .Q(OPER_B[8]), 
        .QN(N169) );
  DFFRX2TF \wtemp_reg[2]  ( .D(N680), .CK(CLK), .RN(RST_N), .Q(OPER_B[2]), 
        .QN(N165) );
  DFFRX2TF \wtemp_reg[10]  ( .D(N672), .CK(CLK), .RN(RST_N), .Q(OPER_B[10]), 
        .QN(N170) );
  DFFRX2TF \wtemp_reg[12]  ( .D(N724), .CK(CLK), .RN(RST_N), .Q(OPER_B[12]), 
        .QN(N185) );
  DFFRX2TF \ytemp_reg[6]  ( .D(N688), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[6]), .QN(N158) );
  DFFRX2TF \xtemp_reg[8]  ( .D(N711), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[12]), .QN(N159) );
  DFFRX2TF \xtemp_reg[0]  ( .D(N719), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[4]), .QN(N163) );
  DFFRX2TF \wtemp_reg[0]  ( .D(N682), .CK(CLK), .RN(RST_N), .Q(OPER_B[0]), 
        .QN(N182) );
  DFFRX2TF \ytemp_reg[1]  ( .D(N693), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[1]), .QN(N168) );
  DFFRX2TF \ytemp_reg[2]  ( .D(N692), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[2]), .QN(N164) );
  DFFRX2TF \ytemp_reg[4]  ( .D(N690), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[4]), .QN(N157) );
  DFFRX2TF \ytemp_reg[8]  ( .D(N686), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[8]), .QN(N148) );
  DFFRX2TF \xtemp_reg[2]  ( .D(N717), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[6]), .QN(N151) );
  DFFRX2TF \ytemp_reg[7]  ( .D(N687), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[7]), .QN(N155) );
  DFFRX2TF \wtemp_reg[1]  ( .D(N681), .CK(CLK), .RN(RST_N), .Q(OPER_B[1]), 
        .QN(N180) );
  DFFRX2TF \ytemp_reg[5]  ( .D(N689), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[5]), .QN(N154) );
  DFFRX2TF \wtemp_reg[4]  ( .D(N678), .CK(CLK), .RN(RST_N), .Q(OPER_B[4]), 
        .QN(N175) );
  DFFRX2TF \wtemp_reg[9]  ( .D(N673), .CK(CLK), .RN(RST_N), .Q(OPER_B[9]), 
        .QN(N186) );
  DFFRX2TF \wtemp_reg[11]  ( .D(N671), .CK(CLK), .RN(RST_N), .Q(OPER_B[11]), 
        .QN(N183) );
  DFFRX1TF \ztemp_reg[0]  ( .D(N669), .CK(CLK), .RN(RST_N), .Q(ZTEMP[0]) );
  DFFRX1TF \wtemp_reg[6]  ( .D(N676), .CK(CLK), .RN(RST_N), .Q(OPER_B[6]) );
  DFFRX1TF \ztemp_reg[8]  ( .D(N661), .CK(CLK), .RN(RST_N), .Q(ZTEMP[8]) );
  DFFRX1TF \ztemp_reg[6]  ( .D(N663), .CK(CLK), .RN(RST_N), .Q(ZTEMP[6]) );
  DFFRX1TF \ztemp_reg[4]  ( .D(N665), .CK(CLK), .RN(RST_N), .Q(ZTEMP[4]) );
  DFFRX1TF \ztemp_reg[2]  ( .D(N667), .CK(CLK), .RN(RST_N), .Q(ZTEMP[2]) );
  DFFRX1TF \ztemp_reg[1]  ( .D(N668), .CK(CLK), .RN(RST_N), .Q(ZTEMP[1]) );
  DFFRX1TF \ztemp_reg[5]  ( .D(N664), .CK(CLK), .RN(RST_N), .Q(ZTEMP[5]) );
  DFFRX1TF \ztemp_reg[3]  ( .D(N666), .CK(CLK), .RN(RST_N), .Q(ZTEMP[3]) );
  DFFRX1TF \ztemp_reg[7]  ( .D(N662), .CK(CLK), .RN(RST_N), .Q(ZTEMP[7]) );
  DFFRX1TF \ztemp_reg[9]  ( .D(N660), .CK(CLK), .RN(RST_N), .Q(ZTEMP[9]) );
  DFFRX1TF \ytemp_reg[3]  ( .D(N691), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[3]), .QN(N736) );
  DFFRX1TF \wtemp_reg[5]  ( .D(N677), .CK(CLK), .RN(RST_N), .Q(OPER_B[5]) );
  DFFRX1TF \wtemp_reg[7]  ( .D(N675), .CK(CLK), .RN(RST_N), .Q(OPER_B[7]) );
  DFFRX1TF \ztemp_reg[10]  ( .D(N659), .CK(CLK), .RN(RST_N), .Q(ZTEMP[10]) );
  DFFRX1TF \ztemp_reg[11]  ( .D(N658), .CK(CLK), .RN(RST_N), .Q(ZTEMP[11]) );
  DFFRX1TF \ztemp_reg[12]  ( .D(N657), .CK(CLK), .RN(RST_N), .Q(ZTEMP[12]) );
  DFFRX1TF \xtemp_reg[12]  ( .D(N723), .CK(CLK), .RN(RST_N), .Q(XTEMP[12]), 
        .QN(N352) );
  DFFRX1TF \ytemp_reg[11]  ( .D(N683), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[2]), .QN(N813) );
  DFFRX1TF \ytemp_reg[12]  ( .D(N706), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[3]), .QN(N648) );
  DFFRX2TF \xtemp_reg[1]  ( .D(N718), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[5]), .QN(N511) );
  DFFRX2TF \xtemp_reg[9]  ( .D(N710), .CK(CLK), .RN(RST_N), .Q(XTEMP[9]), .QN(
        N528) );
  DFFRX2TF \xtemp_reg[7]  ( .D(N712), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[11]), .QN(N461) );
  DFFRX2TF \xtemp_reg[5]  ( .D(N714), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[9]), .QN(N439) );
  DFFRX2TF \xtemp_reg[6]  ( .D(N713), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[10]), .QN(N525) );
  DFFRX2TF \xtemp_reg[4]  ( .D(N715), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[8]), .QN(N520) );
  DFFRX2TF sign_x_reg ( .D(N722), .CK(CLK), .RN(RST_N), .Q(N961), .QN(N74) );
  DFFRX2TF \index_reg[2]  ( .D(N698), .CK(CLK), .RN(RST_N), .Q(\INDEX[2] ) );
  OA21XLTF U3 ( .A0(SUM_AB[12]), .A1(N650), .B0(N127), .Y(N144) );
  NAND2X1TF U4 ( .A(PRE_WORK), .B(N967), .Y(N382) );
  CLKBUFX2TF U5 ( .A(N255), .Y(N188) );
  CLKBUFX2TF U6 ( .A(N188), .Y(N143) );
  AOI32XLTF U7 ( .A0(N822), .A1(N84), .A2(N823), .B0(N637), .B1(N942), .Y(N643) );
  AOI211X2TF U8 ( .A0(N570), .A1(N84), .B0(N594), .C0(N569), .Y(N596) );
  AND2X2TF U9 ( .A(N215), .B(PRE_WORK), .Y(DP_OP_333_124_4748_N57) );
  AOI21X1TF U10 ( .A0(N826), .A1(N926), .B0(N841), .Y(N1) );
  NOR3X1TF U11 ( .A(OPER_A[1]), .B(N929), .C(N826), .Y(N2) );
  OAI32X1TF U12 ( .A0(N180), .A1(OPER_B[0]), .A2(N119), .B0(N930), .B1(N180), 
        .Y(N3) );
  AOI211X1TF U13 ( .A0(OPER_B[2]), .A1(N851), .B0(N2), .C0(N3), .Y(N4) );
  OAI31X1TF U14 ( .A0(N119), .A1(N182), .A2(OPER_B[1]), .B0(N825), .Y(N5) );
  AOI211X1TF U15 ( .A0(C152_DATA4_1), .A1(N117), .B0(N878), .C0(N5), .Y(N6) );
  OAI211X1TF U16 ( .A0(N827), .A1(N1), .B0(N4), .C0(N6), .Y(N681) );
  AOI22X1TF U17 ( .A0(N1007), .A1(ZTEMP[0]), .B0(N110), .B1(DIVISION_HEAD[0]), 
        .Y(N7) );
  AOI32XLTF U18 ( .A0(N1006), .A1(N7), .A2(N1015), .B0(N972), .B1(N7), .Y(N669) );
  AOI32X1TF U19 ( .A0(N119), .A1(N832), .A2(N930), .B0(N182), .B1(N832), .Y(N8) );
  AOI211X1TF U20 ( .A0(C152_DATA4_0), .A1(N117), .B0(N878), .C0(N8), .Y(N9) );
  OAI21X1TF U21 ( .A0(N841), .A1(N926), .B0(OPER_A[0]), .Y(N10) );
  OAI211X1TF U22 ( .A0(N180), .A1(N881), .B0(N9), .C0(N10), .Y(N682) );
  NOR2X1TF U23 ( .A(N928), .B(OPER_A[11]), .Y(N11) );
  XNOR2X1TF U24 ( .A(OPER_A[12]), .B(N11), .Y(N12) );
  AOI22X1TF U25 ( .A0(N12), .A1(N926), .B0(OPER_A[12]), .B1(N841), .Y(N13) );
  OAI21X1TF U26 ( .A0(N136), .A1(N548), .B0(N125), .Y(N14) );
  XNOR2X1TF U27 ( .A(N14), .B(N85), .Y(N15) );
  XNOR2X1TF U28 ( .A(DP_OP_333_124_4748_N1), .B(N15), .Y(N16) );
  NOR2X1TF U29 ( .A(OPER_B[11]), .B(N931), .Y(N17) );
  OAI31X1TF U30 ( .A0(N118), .A1(N17), .A2(OPER_B[12]), .B0(N825), .Y(N18) );
  AOI211X1TF U31 ( .A0(N117), .A1(N16), .B0(N924), .C0(N18), .Y(N19) );
  OAI31X1TF U32 ( .A0(OPER_B[11]), .A1(N931), .A2(N905), .B0(N861), .Y(N20) );
  AOI32X1TF U33 ( .A0(N942), .A1(OPER_B[12]), .A2(N20), .B0(N214), .B1(
        OPER_B[12]), .Y(N21) );
  NAND4BX1TF U34 ( .AN(N821), .B(N13), .C(N19), .D(N21), .Y(N724) );
  OAI21X1TF U35 ( .A0(N306), .A1(N628), .B0(N621), .Y(N22) );
  AOI21X1TF U36 ( .A0(N184), .A1(N22), .B0(N378), .Y(N23) );
  NAND4X1TF U37 ( .A(N124), .B(N617), .C(N624), .D(\INDEX[2] ), .Y(N24) );
  NAND4X1TF U38 ( .A(N356), .B(N23), .C(N804), .D(N24), .Y(N725) );
  CLKINVX1TF U39 ( .A(N831), .Y(N25) );
  AOI211X1TF U40 ( .A0(N826), .A1(N827), .B0(N910), .C0(OPER_A[2]), .Y(N26) );
  AOI31X1TF U41 ( .A0(N916), .A1(N165), .A2(N25), .B0(N26), .Y(N27) );
  OAI31X1TF U42 ( .A0(OPER_A[0]), .A1(OPER_A[1]), .A2(N910), .B0(N830), .Y(N28) );
  AOI22X1TF U43 ( .A0(OPER_B[3]), .A1(N914), .B0(OPER_A[2]), .B1(N28), .Y(N29)
         );
  AOI32X1TF U44 ( .A0(N916), .A1(OPER_B[2]), .A2(N831), .B0(N915), .B1(
        OPER_B[2]), .Y(N30) );
  AOI31X1TF U45 ( .A0(N27), .A1(N29), .A2(N30), .B0(N918), .Y(N31) );
  AND4X1TF U46 ( .A(N961), .B(N109), .C(N176), .D(N217), .Y(N32) );
  OAI2BB2XLTF U47 ( .B0(N165), .B1(N923), .A0N(N117), .A1N(C152_DATA4_2), .Y(
        N33) );
  OR4X1TF U48 ( .A(N875), .B(N31), .C(N32), .D(N33), .Y(N680) );
  NOR3X1TF U49 ( .A(Y_IN[12]), .B(Y_IN[11]), .C(Y_IN[10]), .Y(N34) );
  CLKINVX1TF U50 ( .A(N438), .Y(N35) );
  AOI22X1TF U51 ( .A0(N309), .A1(N35), .B0(N738), .B1(N107), .Y(N36) );
  OAI21X1TF U52 ( .A0(X_IN[4]), .A1(N308), .B0(N98), .Y(N37) );
  OAI22X1TF U53 ( .A0(N738), .A1(N107), .B0(X_IN[6]), .B1(N730), .Y(N38) );
  AOI31X1TF U54 ( .A0(N310), .A1(N36), .A2(N37), .B0(N38), .Y(N39) );
  AOI21X1TF U55 ( .A0(N730), .A1(X_IN[6]), .B0(N39), .Y(N40) );
  OA22X1TF U56 ( .A0(N41), .A1(N40), .B0(N486), .B1(N190), .Y(N42) );
  AO21X1TF U57 ( .A0(N466), .A1(N40), .B0(Y_IN[4]), .Y(N43) );
  AOI22X1TF U58 ( .A0(N486), .A1(N190), .B0(N42), .B1(N43), .Y(N44) );
  AOI2BB2X1TF U59 ( .B0(X_IN[9]), .B1(N44), .A0N(N499), .A1N(N97), .Y(N45) );
  CLKINVX1TF U60 ( .A(N44), .Y(N46) );
  AO21X1TF U61 ( .A0(N498), .A1(N46), .B0(Y_IN[6]), .Y(N47) );
  AOI22X1TF U62 ( .A0(N499), .A1(N97), .B0(N45), .B1(N47), .Y(N48) );
  AOI222XLTF U63 ( .A0(N762), .A1(X_IN[11]), .B0(N762), .B1(N48), .C0(X_IN[11]), .C1(N48), .Y(N49) );
  OAI21X1TF U64 ( .A0(Y_IN[9]), .A1(N299), .B0(N49), .Y(N50) );
  OAI211X1TF U65 ( .A0(X_IN[12]), .A1(N784), .B0(N34), .C0(N50), .Y(N770) );
  CLKINVX1TF U66 ( .A(X_IN[7]), .Y(N41) );
  OAI21X1TF U67 ( .A0(N880), .A1(N929), .B0(N927), .Y(N51) );
  AO21X1TF U68 ( .A0(N879), .A1(N932), .B0(N877), .Y(N52) );
  AOI22X1TF U69 ( .A0(OPER_A[7]), .A1(N51), .B0(OPER_B[7]), .B1(N52), .Y(N53)
         );
  OAI31X1TF U70 ( .A0(N879), .A1(N118), .A2(OPER_B[7]), .B0(N53), .Y(N54) );
  AOI211X1TF U71 ( .A0(C152_DATA4_7), .A1(N116), .B0(N202), .C0(N54), .Y(N55)
         );
  NAND3BX1TF U72 ( .AN(OPER_A[7]), .B(N880), .C(N926), .Y(N56) );
  OAI211X1TF U73 ( .A0(N881), .A1(N169), .B0(N55), .C0(N56), .Y(N675) );
  NOR3X1TF U74 ( .A(N948), .B(N947), .C(N135), .Y(N57) );
  AOI211X1TF U75 ( .A0(N946), .A1(N84), .B0(N966), .C0(N57), .Y(N58) );
  OAI22X1TF U76 ( .A0(N941), .A1(N127), .B0(N940), .B1(N969), .Y(N59) );
  NOR4XLTF U77 ( .A(N945), .B(N943), .C(N944), .D(N59), .Y(N60) );
  MXI2X1TF U78 ( .A(N58), .B(N123), .S0(N60), .Y(N670) );
  OR2X2TF U79 ( .A(N342), .B(N599), .Y(N61) );
  INVX2TF U80 ( .A(N967), .Y(N135) );
  INVX2TF U81 ( .A(N942), .Y(N126) );
  INVX2TF U82 ( .A(N126), .Y(N84) );
  OR3X1TF U83 ( .A(PRE_WORK), .B(N605), .C(N599), .Y(N62) );
  NAND2X2TF U84 ( .A(SIGN_Y), .B(N961), .Y(N968) );
  AOI22XLTF U85 ( .A0(DIVISION_HEAD[10]), .A1(N547), .B0(DIVISION_HEAD[9]), 
        .B1(N784), .Y(N323) );
  INVX2TF U86 ( .A(N123), .Y(N65) );
  NAND2X1TF U87 ( .A(N774), .B(N766), .Y(N391) );
  NAND2XLTF U88 ( .A(N800), .B(SUM_AB[8]), .Y(N420) );
  NAND2X1TF U89 ( .A(N923), .B(N199), .Y(N213) );
  CLKINVX1TF U90 ( .A(SUM_AB[4]), .Y(N385) );
  AO21X1TF U91 ( .A0(N777), .A1(N368), .B0(N823), .Y(N506) );
  CLKINVX2TF U92 ( .A(OPER_A[4]), .Y(N849) );
  CLKINVX1TF U93 ( .A(N854), .Y(N852) );
  AND2X2TF U94 ( .A(ZTEMP[5]), .B(N188), .Y(POUT[5]) );
  AND2X2TF U95 ( .A(ZTEMP[7]), .B(N188), .Y(POUT[7]) );
  AND2X2TF U96 ( .A(ZTEMP[6]), .B(N188), .Y(POUT[6]) );
  CLKBUFX2TF U97 ( .A(ALU_START), .Y(N87) );
  CLKINVX1TF U98 ( .A(N190), .Y(N197) );
  CLKINVX1TF U99 ( .A(N620), .Y(N622) );
  CLKINVX1TF U100 ( .A(Y_IN[6]), .Y(N196) );
  CLKINVX1TF U101 ( .A(X_IN[2]), .Y(N772) );
  AOI211X1TF U102 ( .A0(X_IN[3]), .A1(N747), .B0(N436), .C0(N435), .Y(N437) );
  AOI211X1TF U103 ( .A0(X_IN[5]), .A1(N747), .B0(N455), .C0(N454), .Y(N456) );
  AOI211X1TF U104 ( .A0(Y_IN[7]), .A1(N747), .B0(N788), .C0(N787), .Y(N789) );
  OA21XLTF U105 ( .A0(SUM_AB[12]), .A1(N390), .B0(N127), .Y(N502) );
  CLKINVX2TF U106 ( .A(N858), .Y(N207) );
  AND2X2TF U107 ( .A(N891), .B(N916), .Y(N932) );
  INVX1TF U108 ( .A(N894), .Y(N876) );
  OR2X2TF U109 ( .A(N1007), .B(N135), .Y(N1008) );
  AOI22X1TF U110 ( .A0(X_IN[5]), .A1(N441), .B0(N86), .B1(N105), .Y(N443) );
  OAI31X1TF U111 ( .A0(N279), .A1(X_IN[11]), .A2(N547), .B0(N278), .Y(N280) );
  OAI21X1TF U112 ( .A0(N374), .A1(N747), .B0(N376), .Y(N375) );
  AOI22X1TF U113 ( .A0(X_IN[2]), .A1(N139), .B0(X_IN[3]), .B1(N807), .Y(N786)
         );
  AOI22X1TF U114 ( .A0(X_IN[12]), .A1(N807), .B0(X_IN[11]), .B1(N139), .Y(N432) );
  AOI22X1TF U115 ( .A0(Y_IN[9]), .A1(N802), .B0(X_IN[4]), .B1(N139), .Y(N803)
         );
  AOI22X1TF U116 ( .A0(XTEMP[11]), .A1(N134), .B0(N86), .B1(N441), .Y(N348) );
  AOI21X1TF U117 ( .A0(N642), .A1(N942), .B0(N641), .Y(N645) );
  OAI31X1TF U118 ( .A0(N564), .A1(N565), .A2(N563), .B0(N84), .Y(N581) );
  NAND3XLTF U119 ( .A(N942), .B(N824), .C(N823), .Y(N632) );
  INVX1TF U120 ( .A(N400), .Y(N401) );
  OR2X2TF U121 ( .A(N382), .B(N764), .Y(N801) );
  NAND4XLTF U122 ( .A(N611), .B(N610), .C(N609), .D(N608), .Y(N612) );
  OAI31XLTF U123 ( .A0(N127), .A1(N172), .A2(N631), .B0(N630), .Y(N636) );
  OAI2BB2XLTF U124 ( .B0(N762), .B1(N804), .A0N(Y_IN[6]), .A1N(N802), .Y(N779)
         );
  AOI22X1TF U125 ( .A0(X_IN[2]), .A1(N441), .B0(X_IN[1]), .B1(N802), .Y(N414)
         );
  AOI22X1TF U126 ( .A0(DIVISION_HEAD[2]), .A1(N131), .B0(Y_IN[8]), .B1(N802), 
        .Y(N795) );
  NAND3BXLTF U127 ( .AN(N377), .B(N777), .C(N638), .Y(N361) );
  AOI22X1TF U128 ( .A0(N190), .A1(N802), .B0(Y_IN[7]), .B1(N791), .Y(N755) );
  AOI22X1TF U129 ( .A0(Y_IN[3]), .A1(N802), .B0(DIVISION_REMA[6]), .B1(N131), 
        .Y(N742) );
  AOI22X1TF U130 ( .A0(Y_IN[1]), .A1(N802), .B0(DIVISION_REMA[4]), .B1(N131), 
        .Y(N731) );
  OAI211XLTF U131 ( .A0(N136), .A1(N360), .B0(N969), .C0(N600), .Y(N362) );
  OAI21XLTF U132 ( .A0(N135), .A1(N656), .B0(N120), .Y(C2_Z_0) );
  INVX2TF U133 ( .A(N735), .Y(N103) );
  INVX1TF U134 ( .A(OPER_A[11]), .Y(N925) );
  INVX1TF U135 ( .A(OPER_A[8]), .Y(N884) );
  INVX1TF U136 ( .A(OPER_A[1]), .Y(N827) );
  INVX1TF U137 ( .A(OPER_A[10]), .Y(N909) );
  INVX1TF U138 ( .A(OPER_A[6]), .Y(N868) );
  INVX2TF U139 ( .A(N135), .Y(N85) );
  INVX2TF U140 ( .A(N747), .Y(N101) );
  AOI22X1TF U141 ( .A0(DIVISION_REMA[1]), .A1(N112), .B0(ZTEMP[1]), .B1(N173), 
        .Y(N241) );
  AOI22X1TF U142 ( .A0(DIVISION_HEAD[0]), .A1(N113), .B0(ZTEMP[9]), .B1(N65), 
        .Y(N249) );
  AOI22X1TF U143 ( .A0(DIVISION_REMA[5]), .A1(N113), .B0(ZTEMP[5]), .B1(N173), 
        .Y(N245) );
  AOI22X1TF U144 ( .A0(DIVISION_REMA[0]), .A1(N112), .B0(ZTEMP[0]), .B1(N173), 
        .Y(N240) );
  AOI22X1TF U145 ( .A0(DIVISION_HEAD[2]), .A1(N113), .B0(ZTEMP[11]), .B1(N65), 
        .Y(N251) );
  AOI22X1TF U146 ( .A0(DIVISION_REMA[6]), .A1(N113), .B0(ZTEMP[6]), .B1(N173), 
        .Y(N246) );
  AOI22X1TF U147 ( .A0(DIVISION_HEAD[1]), .A1(N113), .B0(ZTEMP[10]), .B1(N65), 
        .Y(N250) );
  AOI22X1TF U148 ( .A0(DIVISION_REMA[4]), .A1(N113), .B0(ZTEMP[4]), .B1(N173), 
        .Y(N244) );
  AOI22X1TF U149 ( .A0(DIVISION_REMA[7]), .A1(N113), .B0(ZTEMP[7]), .B1(N173), 
        .Y(N247) );
  AOI22X1TF U150 ( .A0(DIVISION_REMA[8]), .A1(N113), .B0(ZTEMP[8]), .B1(N173), 
        .Y(N248) );
  AOI22X1TF U151 ( .A0(DIVISION_REMA[2]), .A1(N112), .B0(ZTEMP[2]), .B1(N173), 
        .Y(N242) );
  AOI22X1TF U152 ( .A0(DIVISION_REMA[3]), .A1(N113), .B0(ZTEMP[3]), .B1(N173), 
        .Y(N243) );
  CLKAND2X2TF U153 ( .A(N646), .B(N639), .Y(N545) );
  AND2X2TF U154 ( .A(N379), .B(N345), .Y(N735) );
  AOI22X1TF U155 ( .A0(DIVISION_HEAD[3]), .A1(N113), .B0(ZTEMP[12]), .B1(N65), 
        .Y(N253) );
  INVX2TF U156 ( .A(N61), .Y(N130) );
  INVX2TF U157 ( .A(N252), .Y(N112) );
  INVX1TF U158 ( .A(N336), .Y(N951) );
  AND2X2TF U159 ( .A(N336), .B(N215), .Y(N942) );
  AND2X2TF U160 ( .A(N345), .B(DP_OP_333_124_4748_N57), .Y(N747) );
  NAND2XLTF U161 ( .A(N215), .B(N946), .Y(N533) );
  INVX2TF U162 ( .A(N340), .Y(N341) );
  AND2X2TF U163 ( .A(N123), .B(N239), .Y(N254) );
  OR2X2TF U164 ( .A(N173), .B(N239), .Y(N252) );
  INVX2TF U165 ( .A(N193), .Y(N107) );
  AND2X2TF U166 ( .A(N216), .B(N87), .Y(N967) );
  INVX2TF U167 ( .A(N191), .Y(N97) );
  AND2X2TF U168 ( .A(N63), .B(N188), .Y(N237) );
  AND2X2TF U169 ( .A(N188), .B(N108), .Y(N236) );
  NAND2XLTF U170 ( .A(DIVISION_HEAD[4]), .B(N256), .Y(N218) );
  INVX1TF U171 ( .A(N256), .Y(N141) );
  AOI22X1TF U172 ( .A0(X_IN[11]), .A1(N547), .B0(X_IN[12]), .B1(N805), .Y(N274) );
  INVX2TF U173 ( .A(Y_IN[7]), .Y(N191) );
  INVX2TF U174 ( .A(X_IN[3]), .Y(N192) );
  INVX2TF U175 ( .A(X_IN[5]), .Y(N193) );
  INVX2TF U176 ( .A(N295), .Y(N86) );
  INVX2TF U177 ( .A(N237), .Y(N88) );
  INVX2TF U178 ( .A(N237), .Y(N89) );
  INVX2TF U179 ( .A(N236), .Y(N93) );
  INVX2TF U180 ( .A(N236), .Y(N94) );
  INVX2TF U181 ( .A(N1015), .Y(N95) );
  INVX2TF U182 ( .A(N1015), .Y(N96) );
  INVX2TF U183 ( .A(N192), .Y(N98) );
  INVX2TF U184 ( .A(N62), .Y(N99) );
  INVX2TF U185 ( .A(N62), .Y(N100) );
  INVX2TF U186 ( .A(N747), .Y(N102) );
  INVX2TF U187 ( .A(N735), .Y(N104) );
  INVX2TF U188 ( .A(N391), .Y(N105) );
  INVX2TF U189 ( .A(N391), .Y(N106) );
  INVX2TF U190 ( .A(N108), .Y(N109) );
  INVX2TF U191 ( .A(N1008), .Y(N110) );
  INVX2TF U192 ( .A(N1008), .Y(N111) );
  INVX2TF U193 ( .A(N252), .Y(N113) );
  INVX2TF U194 ( .A(N254), .Y(N114) );
  INVX2TF U195 ( .A(N254), .Y(N115) );
  INVX2TF U196 ( .A(N213), .Y(N116) );
  INVX2TF U197 ( .A(N213), .Y(N117) );
  INVX2TF U198 ( .A(N932), .Y(N118) );
  INVX2TF U199 ( .A(N932), .Y(N119) );
  INVX2TF U200 ( .A(DP_OP_333_124_4748_N57), .Y(N120) );
  INVX2TF U201 ( .A(DP_OP_333_124_4748_N57), .Y(N125) );
  INVX2TF U202 ( .A(N942), .Y(N127) );
  INVX2TF U203 ( .A(N61), .Y(N131) );
  INVX2TF U204 ( .A(N506), .Y(N132) );
  INVX2TF U205 ( .A(N506), .Y(N133) );
  INVX2TF U206 ( .A(N103), .Y(N134) );
  INVX2TF U207 ( .A(N967), .Y(N136) );
  AOI222X4TF U208 ( .A0(N485), .A1(N160), .B0(N485), .B1(N499), .C0(N160), 
        .C1(N499), .Y(N495) );
  NOR2X2TF U209 ( .A(N333), .B(N952), .Y(N345) );
  NOR2X2TF U210 ( .A(N342), .B(N135), .Y(N379) );
  NOR3X2TF U211 ( .A(N126), .B(N604), .C(N631), .Y(N617) );
  INVX2TF U212 ( .A(N502), .Y(N137) );
  INVX2TF U213 ( .A(N502), .Y(N138) );
  INVX2TF U214 ( .A(N801), .Y(N139) );
  INVX2TF U215 ( .A(N801), .Y(N140) );
  NAND2X2TF U216 ( .A(N123), .B(N763), .Y(N451) );
  AOI21X2TF U217 ( .A0(N84), .A1(N915), .B0(N214), .Y(N930) );
  NAND2X2TF U218 ( .A(N564), .B(N341), .Y(N910) );
  AOI22XLTF U219 ( .A0(X_IN[2]), .A1(N802), .B0(X_IN[3]), .B1(N441), .Y(N421)
         );
  INVX2TF U220 ( .A(N965), .Y(N142) );
  AOI2BB1X2TF U221 ( .A0N(N959), .A1N(N958), .B0(N957), .Y(N1007) );
  OAI21XLTF U222 ( .A0(N600), .A1(N599), .B0(N598), .Y(N601) );
  INVXLTF U223 ( .A(N599), .Y(N566) );
  NOR3BX2TF U224 ( .AN(ALU_TYPE[2]), .B(ALU_TYPE[0]), .C(ALU_TYPE[1]), .Y(N256) );
  NOR3XLTF U225 ( .A(N108), .B(N904), .C(N968), .Y(N821) );
  NAND2X2TF U226 ( .A(N966), .B(N923), .Y(N904) );
  AOI21XLTF U227 ( .A0(N822), .A1(N370), .B0(N369), .Y(N372) );
  AOI21XLTF U228 ( .A0(N824), .A1(N823), .B0(N822), .Y(N828) );
  INVXLTF U229 ( .A(N822), .Y(N373) );
  NOR3BX4TF U230 ( .AN(N381), .B(N378), .C(N134), .Y(N510) );
  AOI21X2TF U231 ( .A0(N767), .A1(N303), .B0(N382), .Y(N378) );
  AOI222X4TF U232 ( .A0(XTEMP[9]), .A1(X_IN[9]), .B0(XTEMP[9]), .B1(N476), 
        .C0(X_IN[9]), .C1(N476), .Y(N485) );
  AOI222X4TF U233 ( .A0(N159), .A1(N486), .B0(N159), .B1(N462), .C0(N486), 
        .C1(N462), .Y(N476) );
  OAI21X2TF U234 ( .A0(N511), .A1(N114), .B0(N241), .Y(OPER_A[1]) );
  NAND2X2TF U235 ( .A(N763), .B(N65), .Y(N558) );
  NOR2X4TF U236 ( .A(N382), .B(N769), .Y(N807) );
  AOI22XLTF U237 ( .A0(DIVISION_HEAD[5]), .A1(N99), .B0(X_IN[7]), .B1(N807), 
        .Y(N384) );
  AOI22XLTF U238 ( .A0(X_IN[10]), .A1(N139), .B0(X_IN[11]), .B1(N807), .Y(N423) );
  NOR4X2TF U239 ( .A(N647), .B(N943), .C(N362), .D(N361), .Y(N641) );
  NOR2X2TF U240 ( .A(N333), .B(N603), .Y(N565) );
  NOR2BX2TF U241 ( .AN(N543), .B(N379), .Y(N628) );
  INVX2TF U242 ( .A(N144), .Y(N145) );
  INVX2TF U243 ( .A(N144), .Y(N146) );
  AOI22X2TF U244 ( .A0(N340), .A1(N338), .B0(N941), .B1(N341), .Y(N916) );
  XNOR2X1TF U245 ( .A(OPER_A[12]), .B(ADD_X_132_1_N2), .Y(N147) );
  CMPR32X2TF U246 ( .A(OPER_A[7]), .B(OPER_B[7]), .C(ADD_X_132_1_N7), .CO(
        ADD_X_132_1_N6), .S(SUM_AB[7]) );
  CMPR32X2TF U247 ( .A(OPER_A[6]), .B(OPER_B[6]), .C(ADD_X_132_1_N8), .CO(
        ADD_X_132_1_N7), .S(SUM_AB[6]) );
  XNOR2X2TF U248 ( .A(N147), .B(OPER_B[12]), .Y(SUM_AB[12]) );
  INVX2TF U249 ( .A(OPER_A[0]), .Y(N826) );
  OAI21X2TF U250 ( .A0(N163), .A1(N114), .B0(N240), .Y(OPER_A[0]) );
  NOR2X1TF U251 ( .A(ALU_TYPE[2]), .B(ALU_TYPE[0]), .Y(N194) );
  AOI222XLTF U252 ( .A0(DIVISION_HEAD[1]), .A1(DIVISION_HEAD[0]), .B0(
        DIVISION_HEAD[1]), .B1(N309), .C0(DIVISION_HEAD[0]), .C1(N308), .Y(
        N311) );
  AOI22X1TF U253 ( .A0(N108), .A1(N171), .B0(POST_WORK), .B1(N63), .Y(N239) );
  NAND2X1TF U254 ( .A(N308), .B(N656), .Y(N310) );
  NOR2X1TF U255 ( .A(SUM_AB[10]), .B(N484), .Y(N497) );
  NAND2X1TF U256 ( .A(N475), .B(N474), .Y(N484) );
  NOR2X1TF U257 ( .A(SUM_AB[8]), .B(N459), .Y(N475) );
  OA22X1TF U258 ( .A0(N769), .A1(N557), .B0(N764), .B1(N765), .Y(N303) );
  INVX2TF U259 ( .A(N923), .Y(N214) );
  OAI21X1TF U260 ( .A0(N947), .A1(N609), .B0(N646), .Y(N957) );
  NOR2X2TF U261 ( .A(N214), .B(N126), .Y(N891) );
  OR2X2TF U262 ( .A(N957), .B(N195), .Y(N923) );
  NOR2X1TF U263 ( .A(\INDEX[2] ), .B(N620), .Y(N306) );
  NAND2X1TF U264 ( .A(N129), .B(N128), .Y(N620) );
  OAI21X1TF U265 ( .A0(DIVISION_HEAD[12]), .A1(N548), .B0(N332), .Y(N947) );
  AOI2BB1X1TF U266 ( .A0N(DIVISION_HEAD[6]), .A1N(N321), .B0(Y_IN[6]), .Y(N319) );
  AOI21X1TF U267 ( .A0(N190), .A1(N511), .B0(N318), .Y(N321) );
  AOI2BB1X1TF U268 ( .A0N(DIVISION_HEAD[4]), .A1N(N317), .B0(Y_IN[4]), .Y(N315) );
  NAND2X1TF U269 ( .A(N906), .B(N891), .Y(N927) );
  AOI2BB1X1TF U270 ( .A0N(N607), .A1N(N337), .B0(N958), .Y(N195) );
  NOR2X1TF U271 ( .A(PRE_WORK), .B(N334), .Y(N336) );
  NAND2X1TF U272 ( .A(N122), .B(N161), .Y(N604) );
  NOR2X1TF U273 ( .A(N124), .B(N627), .Y(N334) );
  NAND2X1TF U274 ( .A(N87), .B(N256), .Y(N599) );
  NAND2X1TF U275 ( .A(N565), .B(N379), .Y(N609) );
  NOR2X1TF U276 ( .A(Y_IN[3]), .B(N648), .Y(N313) );
  NAND2X1TF U277 ( .A(N150), .B(N162), .Y(N333) );
  AOI211X1TF U278 ( .A0(N215), .A1(N607), .B0(N945), .C0(N606), .Y(N610) );
  NAND2X1TF U279 ( .A(N451), .B(N457), .Y(N469) );
  NAND2X2TF U280 ( .A(N546), .B(N381), .Y(N457) );
  CLKBUFX2TF U281 ( .A(N782), .Y(N189) );
  AOI211X1TF U282 ( .A0(Y_IN[11]), .A1(N299), .B0(Y_IN[12]), .C0(N280), .Y(
        N767) );
  NAND2X1TF U283 ( .A(N121), .B(N122), .Y(N952) );
  NAND3X1TF U284 ( .A(N958), .B(N135), .C(N599), .Y(N646) );
  AND2X2TF U285 ( .A(N87), .B(N143), .Y(N215) );
  NAND2X1TF U286 ( .A(N174), .B(N360), .Y(N342) );
  NAND2X1TF U287 ( .A(N124), .B(N306), .Y(N360) );
  NAND2X1TF U288 ( .A(N121), .B(N172), .Y(N603) );
  CLKBUFX2TF U289 ( .A(Y_IN[5]), .Y(N190) );
  AND2X2TF U290 ( .A(N194), .B(ALU_TYPE[1]), .Y(N216) );
  NOR3X1TF U291 ( .A(N605), .B(N604), .C(N777), .Y(N606) );
  OR3X1TF U292 ( .A(N875), .B(N874), .C(N209), .Y(N676) );
  OAI2BB2XLTF U293 ( .B0(N876), .B1(N968), .A0N(C152_DATA4_6), .A1N(N117), .Y(
        N209) );
  OAI2BB2XLTF U294 ( .B0(N873), .B1(N918), .A0N(N214), .A1N(OPER_B[6]), .Y(
        N874) );
  INVX2TF U295 ( .A(N457), .Y(N473) );
  AOI32X1TF U296 ( .A0(N966), .A1(N965), .A2(N964), .B0(N942), .B1(N965), .Y(
        N1015) );
  NAND2X1TF U297 ( .A(N565), .B(DP_OP_333_124_4748_N57), .Y(N390) );
  NAND2X1TF U298 ( .A(N956), .B(DP_OP_333_124_4748_N57), .Y(N650) );
  INVX2TF U299 ( .A(N359), .Y(N763) );
  NAND2X1TF U300 ( .A(N379), .B(N956), .Y(N359) );
  NOR2BX2TF U301 ( .AN(N546), .B(N556), .Y(N814) );
  NOR2X1TF U302 ( .A(N174), .B(N599), .Y(N347) );
  NAND2X1TF U303 ( .A(N891), .B(N864), .Y(N881) );
  NOR2X1TF U304 ( .A(N109), .B(N904), .Y(N894) );
  AOI21X1TF U305 ( .A0(N948), .A1(N963), .B0(N358), .Y(N966) );
  NAND2X1TF U306 ( .A(N150), .B(STEP[3]), .Y(N631) );
  NOR2X2TF U307 ( .A(N333), .B(N604), .Y(N956) );
  NAND2X1TF U308 ( .A(N334), .B(N174), .Y(N339) );
  NOR3BX1TF U309 ( .AN(ALU_TYPE[0]), .B(ALU_TYPE[1]), .C(ALU_TYPE[2]), .Y(N255) );
  AO22X1TF U310 ( .A0(N367), .A1(XTEMP[12]), .B0(N355), .B1(N961), .Y(N722) );
  AOI32X1TF U311 ( .A0(N963), .A1(N356), .A2(N954), .B0(N969), .B1(N356), .Y(
        N357) );
  NAND2X1TF U312 ( .A(N946), .B(DP_OP_333_124_4748_N57), .Y(N634) );
  NAND2X1TF U313 ( .A(N642), .B(N131), .Y(N614) );
  NAND2X1TF U314 ( .A(N117), .B(C152_DATA4_8), .Y(N210) );
  AOI32X1TF U315 ( .A0(N132), .A1(DIVISION_HEAD[4]), .A2(N750), .B0(N469), 
        .B1(DIVISION_HEAD[4]), .Y(N388) );
  OAI22X1TF U316 ( .A0(N528), .A1(N104), .B0(N486), .B1(N102), .Y(N487) );
  INVX2TF U317 ( .A(N1011), .Y(N1006) );
  OAI2BB2XLTF U318 ( .B0(N109), .B1(N968), .A0N(N968), .A1N(N109), .Y(N970) );
  NOR2X2TF U319 ( .A(N763), .B(N189), .Y(N761) );
  INVX2TF U320 ( .A(N130), .Y(N777) );
  OAI211X1TF U321 ( .A0(N956), .A1(N342), .B0(N566), .C0(N600), .Y(N343) );
  NAND2X1TF U322 ( .A(N646), .B(N101), .Y(N944) );
  NAND2X1TF U323 ( .A(N345), .B(N130), .Y(N543) );
  NOR2X1TF U324 ( .A(N952), .B(N631), .Y(N563) );
  NOR2X1TF U325 ( .A(N604), .B(N950), .Y(N564) );
  NAND2X1TF U326 ( .A(STEP[2]), .B(N162), .Y(N950) );
  INVX2TF U327 ( .A(N215), .Y(N958) );
  OAI32X1TF U328 ( .A0(N649), .A1(N176), .A2(N944), .B0(N648), .B1(N650), .Y(
        N694) );
  OAI21X1TF U329 ( .A0(N174), .A1(N647), .B0(N646), .Y(N695) );
  AOI22X1TF U330 ( .A0(N542), .A1(N108), .B0(N541), .B1(N540), .Y(N707) );
  INVX2TF U331 ( .A(N542), .Y(N540) );
  OAI31X1TF U332 ( .A0(N539), .A1(N538), .A2(N537), .B0(N536), .Y(N541) );
  AOI211X1TF U333 ( .A0(N535), .A1(XTEMP[12]), .B0(N534), .C0(N533), .Y(N536)
         );
  OAI31X1TF U334 ( .A0(DIVISION_HEAD[1]), .A1(N532), .A2(N160), .B0(N531), .Y(
        N535) );
  AOI22X1TF U335 ( .A0(N530), .A1(N529), .B0(XTEMP[11]), .B1(N813), .Y(N531)
         );
  OAI22X1TF U336 ( .A0(DIVISION_HEAD[0]), .A1(N528), .B0(DIVISION_REMA[8]), 
        .B1(N159), .Y(N529) );
  INVX2TF U337 ( .A(N538), .Y(N530) );
  NOR2X1TF U338 ( .A(XTEMP[11]), .B(N813), .Y(N532) );
  OAI22X1TF U339 ( .A0(DIVISION_HEAD[12]), .A1(N148), .B0(XTEMP[12]), .B1(N648), .Y(N537) );
  OAI21X1TF U340 ( .A0(XTEMP[11]), .A1(N813), .B0(N527), .Y(N538) );
  AOI22X1TF U341 ( .A0(DIVISION_HEAD[0]), .A1(N528), .B0(DIVISION_HEAD[1]), 
        .B1(N160), .Y(N527) );
  AOI21X1TF U342 ( .A0(DIVISION_HEAD[11]), .A1(N155), .B0(N526), .Y(N539) );
  AOI211X1TF U343 ( .A0(DIVISION_REMA[6]), .A1(N525), .B0(N524), .C0(N523), 
        .Y(N526) );
  NOR2X1TF U344 ( .A(DIVISION_HEAD[11]), .B(N155), .Y(N523) );
  AOI21X1TF U345 ( .A0(DIVISION_HEAD[9]), .A1(N154), .B0(N521), .Y(N522) );
  AOI211X1TF U346 ( .A0(DIVISION_REMA[4]), .A1(N520), .B0(N519), .C0(N518), 
        .Y(N521) );
  NOR2X1TF U347 ( .A(DIVISION_HEAD[9]), .B(N154), .Y(N518) );
  AOI21X1TF U348 ( .A0(DIVISION_HEAD[7]), .A1(N736), .B0(N516), .Y(N517) );
  AOI211X1TF U349 ( .A0(N515), .A1(DIVISION_REMA[2]), .B0(N514), .C0(N513), 
        .Y(N516) );
  NOR2X1TF U350 ( .A(DIVISION_HEAD[7]), .B(N736), .Y(N514) );
  OAI21X1TF U351 ( .A0(DIVISION_HEAD[5]), .A1(N168), .B0(N512), .Y(N515) );
  OAI211X1TF U352 ( .A0(DIVISION_REMA[1]), .A1(N511), .B0(DIVISION_REMA[0]), 
        .C0(N163), .Y(N512) );
  OAI21X1TF U353 ( .A0(N376), .A1(N171), .B0(N375), .Y(N720) );
  OAI22X1TF U354 ( .A0(N127), .A1(N373), .B0(N764), .B1(N639), .Y(N374) );
  OAI211X1TF U355 ( .A0(N368), .A1(N823), .B0(N611), .C0(N639), .Y(N369) );
  OAI21X1TF U356 ( .A0(N596), .A1(N585), .B0(N584), .Y(N702) );
  AOI31X1TF U357 ( .A0(N583), .A1(N588), .A2(N590), .B0(N582), .Y(N585) );
  OAI22X1TF U358 ( .A0(N128), .A1(N581), .B0(N592), .B1(N588), .Y(N582) );
  AOI22X1TF U359 ( .A0(N596), .A1(N92), .B0(N580), .B1(N579), .Y(N703) );
  AOI211X1TF U360 ( .A0(N594), .A1(N166), .B0(N578), .C0(N791), .Y(N580) );
  AOI21X1TF U361 ( .A0(N577), .A1(N777), .B0(N178), .Y(N578) );
  OAI21X1TF U362 ( .A0(N128), .A1(N619), .B0(N618), .Y(N699) );
  AOI31X1TF U363 ( .A0(N617), .A1(N620), .A2(N616), .B0(N615), .Y(N618) );
  OAI32X1TF U364 ( .A0(N628), .A1(N629), .A2(N620), .B0(N616), .B1(N628), .Y(
        N615) );
  OAI21X1TF U365 ( .A0(N129), .A1(N619), .B0(N305), .Y(N726) );
  OAI21X1TF U366 ( .A0(N304), .A1(N378), .B0(N619), .Y(N305) );
  AOI32X1TF U367 ( .A0(N628), .A1(N634), .A2(N371), .B0(N166), .B1(N634), .Y(
        N304) );
  OAI31X1TF U368 ( .A0(N629), .A1(N628), .A2(N627), .B0(N626), .Y(N698) );
  AOI22X1TF U369 ( .A0(\INDEX[2] ), .A1(N625), .B0(N624), .B1(N623), .Y(N626)
         );
  OAI21X1TF U370 ( .A0(N622), .A1(N628), .B0(N621), .Y(N625) );
  OAI211X1TF U371 ( .A0(N127), .A1(N364), .B0(N644), .C0(N363), .Y(N721) );
  AOI22X1TF U372 ( .A0(STEP[3]), .A1(N641), .B0(N370), .B1(N573), .Y(N363) );
  NOR2X1TF U373 ( .A(N629), .B(N623), .Y(N621) );
  AOI21X1TF U374 ( .A0(\INDEX[2] ), .A1(N624), .B0(N371), .Y(N623) );
  INVX2TF U375 ( .A(N619), .Y(N629) );
  INVX2TF U376 ( .A(N616), .Y(N624) );
  OAI211X1TF U377 ( .A0(N177), .A1(N614), .B0(N630), .C0(N613), .Y(N700) );
  AOI21X1TF U378 ( .A0(N641), .A1(N161), .B0(N612), .Y(N613) );
  NOR3X1TF U379 ( .A(STEP[3]), .B(N127), .C(N603), .Y(N945) );
  AOI211X1TF U380 ( .A0(N824), .A1(N370), .B0(N367), .C0(N366), .Y(N611) );
  AOI21X1TF U381 ( .A0(N380), .A1(N365), .B0(N777), .Y(N366) );
  NOR2X1TF U382 ( .A(N126), .B(N823), .Y(N370) );
  OAI22X1TF U383 ( .A0(N90), .A1(N597), .B0(N596), .B1(N595), .Y(N701) );
  AOI21X1TF U384 ( .A0(\INDEX[2] ), .A1(N594), .B0(N593), .Y(N595) );
  OAI22X1TF U385 ( .A0(N592), .A1(N591), .B0(N590), .B1(N589), .Y(N593) );
  INVX2TF U386 ( .A(N587), .Y(N592) );
  AOI21X1TF U387 ( .A0(N588), .A1(N587), .B0(N586), .Y(N597) );
  OAI211X1TF U388 ( .A0(N645), .A1(N150), .B0(N644), .C0(N643), .Y(N696) );
  NOR2X1TF U389 ( .A(N649), .B(N357), .Y(N644) );
  OAI21X1TF U390 ( .A0(N345), .A1(N257), .B0(N84), .Y(N356) );
  INVX2TF U391 ( .A(N650), .Y(N649) );
  OAI22X1TF U392 ( .A0(N172), .A1(N950), .B0(N823), .B1(N963), .Y(N637) );
  AOI211X1TF U393 ( .A0(N641), .A1(N172), .B0(N636), .C0(N635), .Y(N640) );
  INVX2TF U394 ( .A(N258), .Y(N633) );
  AOI31X1TF U395 ( .A0(N952), .A1(N365), .A2(N380), .B0(N777), .Y(N258) );
  AOI21X1TF U396 ( .A0(N967), .A1(N602), .B0(N601), .Y(N630) );
  OAI22X1TF U397 ( .A0(N596), .A1(N576), .B0(N575), .B1(N187), .Y(N704) );
  AOI21X1TF U398 ( .A0(N591), .A1(N587), .B0(N586), .Y(N575) );
  OAI21X1TF U399 ( .A0(N90), .A1(N590), .B0(N583), .Y(N589) );
  INVX2TF U400 ( .A(N614), .Y(N583) );
  INVX2TF U401 ( .A(N596), .Y(N579) );
  OAI31X1TF U402 ( .A0(N605), .A1(N604), .A2(N777), .B0(N577), .Y(N587) );
  OAI32X1TF U403 ( .A0(N574), .A1(N824), .A2(N573), .B0(N942), .B1(N574), .Y(
        N577) );
  INVX2TF U404 ( .A(N572), .Y(N574) );
  AOI21X1TF U405 ( .A0(N594), .A1(N184), .B0(N571), .Y(N576) );
  AOI32X1TF U406 ( .A0(N565), .A1(N131), .A2(N177), .B0(N956), .B1(N130), .Y(
        N567) );
  AOI31X1TF U407 ( .A0(N84), .A1(N824), .A2(N823), .B0(N944), .Y(N568) );
  INVX2TF U408 ( .A(N581), .Y(N594) );
  AOI22X1TF U409 ( .A0(N890), .A1(N891), .B0(N214), .B1(OPER_B[8]), .Y(N211)
         );
  OAI21X1TF U410 ( .A0(N889), .A1(N169), .B0(N888), .Y(N890) );
  AOI211X1TF U411 ( .A0(N914), .A1(OPER_B[9]), .B0(N887), .C0(N886), .Y(N888)
         );
  OAI32X1TF U412 ( .A0(OPER_A[8]), .A1(N885), .A2(N910), .B0(N884), .B1(N883), 
        .Y(N886) );
  AOI21X1TF U413 ( .A0(N907), .A1(N885), .B0(N906), .Y(N883) );
  NOR3X1TF U414 ( .A(N905), .B(OPER_B[8]), .C(N882), .Y(N887) );
  AOI21X1TF U415 ( .A0(N882), .A1(N916), .B0(N915), .Y(N889) );
  OAI21X1TF U416 ( .A0(N447), .A1(N446), .B0(N457), .Y(N448) );
  AOI22X1TF U417 ( .A0(DIVISION_HEAD[11]), .A1(N100), .B0(X_IN[12]), .B1(N140), 
        .Y(N442) );
  AOI22X1TF U418 ( .A0(SUM_AB[6]), .A1(N137), .B0(N491), .B1(N988), .Y(N444)
         );
  OAI22X1TF U419 ( .A0(N439), .A1(N104), .B0(N438), .B1(N102), .Y(N447) );
  OAI211X1TF U420 ( .A0(N1006), .A1(N993), .B0(N992), .C0(N991), .Y(N662) );
  AOI22X1TF U421 ( .A0(DIVISION_HEAD[7]), .A1(N110), .B0(ZTEMP[7]), .B1(N142), 
        .Y(N992) );
  OAI211X1TF U422 ( .A0(N1006), .A1(N981), .B0(N980), .C0(N979), .Y(N666) );
  AOI22X1TF U423 ( .A0(DIVISION_HEAD[3]), .A1(N110), .B0(ZTEMP[3]), .B1(N1007), 
        .Y(N980) );
  OAI211X1TF U424 ( .A0(N1006), .A1(N987), .B0(N986), .C0(N985), .Y(N664) );
  AOI22X1TF U425 ( .A0(DIVISION_HEAD[5]), .A1(N110), .B0(ZTEMP[5]), .B1(N142), 
        .Y(N986) );
  AOI22X1TF U426 ( .A0(SUM_AB[4]), .A1(N95), .B0(N982), .B1(N1011), .Y(N983)
         );
  AOI22X1TF U427 ( .A0(DIVISION_HEAD[4]), .A1(N111), .B0(ZTEMP[4]), .B1(N142), 
        .Y(N984) );
  AOI22X1TF U428 ( .A0(SUM_AB[8]), .A1(N95), .B0(N994), .B1(N1011), .Y(N995)
         );
  AOI22X1TF U429 ( .A0(DIVISION_HEAD[8]), .A1(N111), .B0(ZTEMP[8]), .B1(N142), 
        .Y(N996) );
  AOI22X1TF U430 ( .A0(SUM_AB[6]), .A1(N95), .B0(N988), .B1(N1011), .Y(N989)
         );
  AOI22X1TF U431 ( .A0(DIVISION_HEAD[6]), .A1(N111), .B0(ZTEMP[6]), .B1(N142), 
        .Y(N990) );
  AOI22X1TF U432 ( .A0(SUM_AB[1]), .A1(N95), .B0(N973), .B1(N1011), .Y(N974)
         );
  AOI22X1TF U433 ( .A0(DIVISION_HEAD[1]), .A1(N111), .B0(ZTEMP[1]), .B1(N142), 
        .Y(N975) );
  AOI22X1TF U434 ( .A0(SUM_AB[2]), .A1(N95), .B0(N976), .B1(N1011), .Y(N977)
         );
  AOI22X1TF U435 ( .A0(DIVISION_HEAD[2]), .A1(N111), .B0(ZTEMP[2]), .B1(N142), 
        .Y(N978) );
  OAI211X1TF U436 ( .A0(N1006), .A1(N999), .B0(N998), .C0(N997), .Y(N660) );
  AOI22X1TF U437 ( .A0(DIVISION_HEAD[9]), .A1(N110), .B0(ZTEMP[9]), .B1(N1007), 
        .Y(N998) );
  AOI211X1TF U438 ( .A0(N214), .A1(OPER_B[10]), .B0(N921), .C0(N922), .Y(N212)
         );
  AOI21X1TF U439 ( .A0(N971), .A1(N968), .B0(N904), .Y(N922) );
  AOI21X1TF U440 ( .A0(N920), .A1(N919), .B0(N918), .Y(N921) );
  AOI32X1TF U441 ( .A0(N917), .A1(OPER_B[10]), .A2(N916), .B0(N915), .B1(
        OPER_B[10]), .Y(N919) );
  AOI211X1TF U442 ( .A0(N914), .A1(OPER_B[11]), .B0(N913), .C0(N912), .Y(N920)
         );
  OAI32X1TF U443 ( .A0(OPER_A[10]), .A1(N911), .A2(N910), .B0(N909), .B1(N908), 
        .Y(N912) );
  AOI21X1TF U444 ( .A0(N907), .A1(N911), .B0(N906), .Y(N908) );
  NOR3X1TF U445 ( .A(N905), .B(OPER_B[10]), .C(N917), .Y(N913) );
  OAI22X1TF U446 ( .A0(N473), .A1(N472), .B0(N471), .B1(N159), .Y(N711) );
  AOI211X1TF U447 ( .A0(N994), .A1(N491), .B0(N468), .C0(N467), .Y(N472) );
  OAI211X1TF U448 ( .A0(N466), .A1(N608), .B0(N465), .C0(N464), .Y(N467) );
  AOI22X1TF U449 ( .A0(XTEMP[9]), .A1(N100), .B0(N800), .B1(SUM_AB[12]), .Y(
        N464) );
  NOR2X1TF U450 ( .A(DIVISION_HEAD[12]), .B(N470), .Y(N463) );
  AOI22X1TF U451 ( .A0(X_IN[8]), .A1(N462), .B0(INTADD_0_N1), .B1(N486), .Y(
        N470) );
  OAI22X1TF U452 ( .A0(N461), .A1(N104), .B0(N460), .B1(N102), .Y(N468) );
  AOI211X1TF U453 ( .A0(OPER_B[6]), .A1(N872), .B0(N871), .C0(N870), .Y(N873)
         );
  OAI32X1TF U454 ( .A0(OPER_A[6]), .A1(N869), .A2(N910), .B0(N868), .B1(N867), 
        .Y(N870) );
  AOI21X1TF U455 ( .A0(N907), .A1(N869), .B0(N906), .Y(N867) );
  INVX2TF U456 ( .A(N910), .Y(N907) );
  OAI31X1TF U457 ( .A0(N905), .A1(OPER_B[6]), .A2(N866), .B0(N865), .Y(N871)
         );
  AOI21X1TF U458 ( .A0(OPER_B[7]), .A1(N864), .B0(N863), .Y(N865) );
  OAI21X1TF U459 ( .A0(N905), .A1(N862), .B0(N861), .Y(N872) );
  AOI32X1TF U460 ( .A0(N427), .A1(N457), .A2(N426), .B0(N473), .B1(N520), .Y(
        N715) );
  AOI211X1TF U461 ( .A0(N491), .A1(N982), .B0(N425), .C0(N424), .Y(N426) );
  AOI22X1TF U462 ( .A0(DIVISION_HEAD[9]), .A1(N99), .B0(X_IN[9]), .B1(N106), 
        .Y(N422) );
  OAI22X1TF U463 ( .A0(N152), .A1(N104), .B0(N520), .B1(N451), .Y(N425) );
  AOI32X1TF U464 ( .A0(N408), .A1(N457), .A2(N407), .B0(N473), .B1(N151), .Y(
        N717) );
  AOI211X1TF U465 ( .A0(DIVISION_HEAD[7]), .A1(N100), .B0(N406), .C0(N405), 
        .Y(N407) );
  OAI211X1TF U466 ( .A0(N102), .A1(N750), .B0(N404), .C0(N403), .Y(N405) );
  AOI21X1TF U467 ( .A0(N491), .A1(N976), .B0(N402), .Y(N403) );
  OAI22X1TF U468 ( .A0(N511), .A1(N103), .B0(N151), .B1(N451), .Y(N402) );
  AOI22X1TF U469 ( .A0(X_IN[1]), .A1(N441), .B0(N800), .B1(SUM_AB[6]), .Y(N404) );
  OAI21X1TF U470 ( .A0(N498), .A1(N749), .B0(N399), .Y(N406) );
  AOI22X1TF U471 ( .A0(X_IN[8]), .A1(N140), .B0(X_IN[7]), .B1(N106), .Y(N399)
         );
  AOI32X1TF U472 ( .A0(N389), .A1(N388), .A2(N387), .B0(N473), .B1(N388), .Y(
        N719) );
  OAI211X1TF U473 ( .A0(N385), .A1(N558), .B0(N384), .C0(N383), .Y(N386) );
  AOI22X1TF U474 ( .A0(X_IN[6]), .A1(N140), .B0(X_IN[5]), .B1(N106), .Y(N383)
         );
  AOI22X1TF U475 ( .A0(DIVISION_HEAD[3]), .A1(N735), .B0(SUM_AB[0]), .B1(N377), 
        .Y(N389) );
  AOI32X1TF U476 ( .A0(N398), .A1(N457), .A2(N397), .B0(N473), .B1(N511), .Y(
        N718) );
  AOI211X1TF U477 ( .A0(N491), .A1(N973), .B0(N396), .C0(N395), .Y(N397) );
  OAI211X1TF U478 ( .A0(N558), .A1(N428), .B0(N394), .C0(N393), .Y(N395) );
  AOI21X1TF U479 ( .A0(DIVISION_HEAD[4]), .A1(N735), .B0(N392), .Y(N393) );
  OAI22X1TF U480 ( .A0(N511), .A1(N451), .B0(N750), .B1(N608), .Y(N392) );
  AOI22X1TF U481 ( .A0(DIVISION_HEAD[6]), .A1(N100), .B0(X_IN[7]), .B1(N139), 
        .Y(N394) );
  OAI22X1TF U482 ( .A0(N460), .A1(N391), .B0(N486), .B1(N749), .Y(N396) );
  AOI32X1TF U483 ( .A0(N458), .A1(N457), .A2(N456), .B0(N473), .B1(N461), .Y(
        N712) );
  OAI211X1TF U484 ( .A0(N504), .A1(N993), .B0(N453), .C0(N452), .Y(N454) );
  AOI22X1TF U485 ( .A0(DIVISION_HEAD[12]), .A1(N99), .B0(X_IN[12]), .B1(N105), 
        .Y(N452) );
  AOI22X1TF U486 ( .A0(DIVISION_HEAD[11]), .A1(N806), .B0(DIVISION_HEAD[10]), 
        .B1(N134), .Y(N453) );
  OAI22X1TF U487 ( .A0(N460), .A1(N608), .B0(N558), .B1(N496), .Y(N455) );
  OAI22X1TF U488 ( .A0(N510), .A1(N483), .B0(N482), .B1(N528), .Y(N710) );
  AOI211X1TF U489 ( .A0(SUM_AB[9]), .A1(N138), .B0(N480), .C0(N479), .Y(N483)
         );
  OAI211X1TF U490 ( .A0(N999), .A1(N504), .B0(N478), .C0(N477), .Y(N479) );
  AOI22X1TF U491 ( .A0(XTEMP[10]), .A1(N100), .B0(X_IN[7]), .B1(N802), .Y(N478) );
  OAI22X1TF U492 ( .A0(N159), .A1(N104), .B0(N486), .B1(N608), .Y(N480) );
  AOI22X1TF U493 ( .A0(N189), .A1(N148), .B0(N781), .B1(N780), .Y(N686) );
  AOI211X1TF U494 ( .A0(DIVISION_REMA[7]), .A1(N735), .B0(N779), .C0(N778), 
        .Y(N781) );
  OAI211X1TF U495 ( .A0(N156), .A1(N777), .B0(N776), .C0(N775), .Y(N778) );
  AOI22X1TF U496 ( .A0(N774), .A1(N773), .B0(N994), .B1(N797), .Y(N775) );
  AOI21X1TF U497 ( .A0(SUM_AB[8]), .A1(N459), .B0(N475), .Y(N994) );
  AOI32X1TF U498 ( .A0(N772), .A1(N771), .A2(N770), .B0(N769), .B1(N771), .Y(
        N773) );
  OAI32X1TF U499 ( .A0(N768), .A1(N767), .A2(X_IN[0]), .B0(N766), .B1(N768), 
        .Y(N771) );
  AOI22X1TF U500 ( .A0(DIVISION_REMA[8]), .A1(N763), .B0(SUM_AB[8]), .B1(N145), 
        .Y(N776) );
  AOI22X1TF U501 ( .A0(SUM_AB[10]), .A1(N96), .B0(N1000), .B1(N1011), .Y(N1001) );
  AOI22X1TF U502 ( .A0(DIVISION_HEAD[10]), .A1(N111), .B0(ZTEMP[10]), .B1(N142), .Y(N1002) );
  AOI22X1TF U503 ( .A0(N473), .A1(N439), .B0(N437), .B1(N457), .Y(N714) );
  AOI21X1TF U504 ( .A0(DIVISION_HEAD[8]), .A1(N134), .B0(N430), .Y(N431) );
  OAI22X1TF U505 ( .A0(N439), .A1(N451), .B0(N504), .B1(N987), .Y(N430) );
  AOI22X1TF U506 ( .A0(DIVISION_HEAD[10]), .A1(N99), .B0(X_IN[10]), .B1(N105), 
        .Y(N433) );
  OAI22X1TF U507 ( .A0(N438), .A1(N608), .B0(N558), .B1(N474), .Y(N436) );
  AOI32X1TF U508 ( .A0(N799), .A1(N816), .A2(N798), .B0(N814), .B1(N149), .Y(
        N684) );
  AOI21X1TF U509 ( .A0(N797), .A1(N1000), .B0(N796), .Y(N798) );
  AOI22X1TF U510 ( .A0(X_IN[2]), .A1(N106), .B0(X_IN[4]), .B1(N807), .Y(N792)
         );
  AOI22X1TF U511 ( .A0(DIVISION_HEAD[0]), .A1(N134), .B0(DIVISION_HEAD[1]), 
        .B1(N806), .Y(N793) );
  AOI22X1TF U512 ( .A0(Y_IN[10]), .A1(N791), .B0(X_IN[3]), .B1(N140), .Y(N794)
         );
  AOI22X1TF U513 ( .A0(N800), .A1(SUM_AB[1]), .B0(SUM_AB[10]), .B1(N146), .Y(
        N799) );
  OAI22X1TF U514 ( .A0(N510), .A1(N494), .B0(N493), .B1(N160), .Y(N709) );
  AOI21X1TF U515 ( .A0(N491), .A1(N1000), .B0(N490), .Y(N494) );
  OAI211X1TF U516 ( .A0(N498), .A1(N608), .B0(N489), .C0(N488), .Y(N490) );
  AOI22X1TF U517 ( .A0(XTEMP[11]), .A1(N100), .B0(SUM_AB[10]), .B1(N137), .Y(
        N489) );
  AOI21X1TF U518 ( .A0(SUM_AB[10]), .A1(N484), .B0(N497), .Y(N1000) );
  AOI32X1TF U519 ( .A0(N418), .A1(N457), .A2(N417), .B0(N473), .B1(N152), .Y(
        N716) );
  AOI211X1TF U520 ( .A0(DIVISION_HEAD[8]), .A1(N100), .B0(N416), .C0(N415), 
        .Y(N417) );
  OAI211X1TF U521 ( .A0(N558), .A1(N449), .B0(N414), .C0(N413), .Y(N415) );
  AOI21X1TF U522 ( .A0(DIVISION_HEAD[6]), .A1(N735), .B0(N412), .Y(N413) );
  OAI22X1TF U523 ( .A0(N152), .A1(N451), .B0(N504), .B1(N981), .Y(N412) );
  OAI21X1TF U524 ( .A0(N499), .A1(N749), .B0(N409), .Y(N416) );
  AOI22X1TF U525 ( .A0(X_IN[8]), .A1(N106), .B0(X_IN[9]), .B1(N140), .Y(N409)
         );
  OAI211X1TF U526 ( .A0(N1006), .A1(N1005), .B0(N1004), .C0(N1003), .Y(N658)
         );
  AOI22X1TF U527 ( .A0(DIVISION_HEAD[11]), .A1(N111), .B0(ZTEMP[11]), .B1(N142), .Y(N1004) );
  OAI21X1TF U528 ( .A0(N761), .A1(N177), .B0(N562), .Y(N705) );
  OAI22X1TF U529 ( .A0(N561), .A1(N560), .B0(N763), .B1(N780), .Y(N562) );
  AOI22X1TF U530 ( .A0(Y_IN[0]), .A1(N791), .B0(DIVISION_REMA[1]), .B1(N130), 
        .Y(N559) );
  AOI21X1TF U531 ( .A0(N127), .A1(N650), .B0(N972), .Y(N561) );
  INVX2TF U532 ( .A(SUM_AB[0]), .Y(N972) );
  OAI22X1TF U533 ( .A0(N189), .A1(N654), .B0(N761), .B1(N168), .Y(N693) );
  AOI21X1TF U534 ( .A0(SUM_AB[1]), .A1(N146), .B0(N653), .Y(N654) );
  AOI22X1TF U535 ( .A0(DIVISION_REMA[0]), .A1(N735), .B0(N797), .B1(N973), .Y(
        N651) );
  AOI21X1TF U536 ( .A0(SUM_AB[1]), .A1(SUM_AB[0]), .B0(N400), .Y(N973) );
  AOI22X1TF U537 ( .A0(Y_IN[1]), .A1(N791), .B0(DIVISION_REMA[2]), .B1(N131), 
        .Y(N652) );
  OAI211X1TF U538 ( .A0(N1015), .A1(N1014), .B0(N1013), .C0(N1012), .Y(N657)
         );
  AOI32X1TF U539 ( .A0(N1014), .A1(N1011), .A2(N1010), .B0(N1009), .B1(N1011), 
        .Y(N1012) );
  AOI211X4TF U540 ( .A0(N971), .A1(N970), .B0(N969), .C0(N1007), .Y(N1011) );
  INVX2TF U541 ( .A(N966), .Y(N969) );
  AOI22X1TF U542 ( .A0(DIVISION_HEAD[12]), .A1(N111), .B0(ZTEMP[12]), .B1(
        N1007), .Y(N1013) );
  OAI31X1TF U543 ( .A0(N963), .A1(N109), .A2(N968), .B0(N962), .Y(N964) );
  AOI31X1TF U544 ( .A0(N176), .A1(N109), .A2(N961), .B0(N960), .Y(N962) );
  INVX2TF U545 ( .A(N1007), .Y(N965) );
  AOI31X1TF U546 ( .A0(N956), .A1(N955), .A2(N954), .B0(N953), .Y(N959) );
  OAI31X1TF U547 ( .A0(N952), .A1(N951), .A2(N950), .B0(N949), .Y(N953) );
  OAI22X1TF U548 ( .A0(N189), .A1(N729), .B0(N761), .B1(N164), .Y(N692) );
  AOI211X1TF U549 ( .A0(SUM_AB[2]), .A1(N146), .B0(N728), .C0(N727), .Y(N729)
         );
  OAI211X1TF U550 ( .A0(N656), .A1(N102), .B0(N757), .C0(N655), .Y(N727) );
  AOI22X1TF U551 ( .A0(DIVISION_REMA[3]), .A1(N131), .B0(N797), .B1(N976), .Y(
        N655) );
  AOI21X1TF U552 ( .A0(SUM_AB[2]), .A1(N401), .B0(N411), .Y(N976) );
  NOR2X1TF U553 ( .A(SUM_AB[0]), .B(SUM_AB[1]), .Y(N400) );
  OAI22X1TF U554 ( .A0(N738), .A1(N804), .B0(N168), .B1(N104), .Y(N728) );
  OAI22X1TF U555 ( .A0(N189), .A1(N753), .B0(N761), .B1(N158), .Y(N688) );
  AOI211X1TF U556 ( .A0(N988), .A1(N797), .B0(N752), .C0(N751), .Y(N753) );
  OAI211X1TF U557 ( .A0(N750), .A1(N749), .B0(N757), .C0(N748), .Y(N751) );
  AOI22X1TF U558 ( .A0(DIVISION_REMA[7]), .A1(N130), .B0(SUM_AB[6]), .B1(N145), 
        .Y(N748) );
  INVX2TF U559 ( .A(N807), .Y(N749) );
  OAI21X1TF U560 ( .A0(N198), .A1(N102), .B0(N746), .Y(N752) );
  AOI22X1TF U561 ( .A0(Y_IN[6]), .A1(N791), .B0(DIVISION_REMA[5]), .B1(N735), 
        .Y(N746) );
  AOI21X1TF U562 ( .A0(SUM_AB[6]), .A1(N440), .B0(N450), .Y(N988) );
  OAI22X1TF U563 ( .A0(N189), .A1(N741), .B0(N761), .B1(N157), .Y(N690) );
  AOI211X1TF U564 ( .A0(SUM_AB[4]), .A1(N146), .B0(N740), .C0(N739), .Y(N741)
         );
  OAI211X1TF U565 ( .A0(N738), .A1(N102), .B0(N757), .C0(N737), .Y(N739) );
  AOI22X1TF U566 ( .A0(DIVISION_REMA[5]), .A1(N131), .B0(N797), .B1(N982), .Y(
        N737) );
  AOI21X1TF U567 ( .A0(SUM_AB[4]), .A1(N419), .B0(N429), .Y(N982) );
  OAI22X1TF U568 ( .A0(N198), .A1(N804), .B0(N736), .B1(N104), .Y(N740) );
  INVX2TF U569 ( .A(N916), .Y(N905) );
  OAI22X1TF U570 ( .A0(N510), .A1(N509), .B0(N508), .B1(N153), .Y(N708) );
  OAI21X1TF U571 ( .A0(N504), .A1(N1005), .B0(N503), .Y(N505) );
  AOI211X1TF U572 ( .A0(SUM_AB[11]), .A1(N137), .B0(N501), .C0(N500), .Y(N503)
         );
  OAI22X1TF U573 ( .A0(N160), .A1(N103), .B0(N498), .B1(N101), .Y(N501) );
  INVX2TF U574 ( .A(N491), .Y(N504) );
  OAI21X1TF U575 ( .A0(N761), .A1(N155), .B0(N760), .Y(N687) );
  OAI21X1TF U576 ( .A0(N759), .A1(N758), .B0(N780), .Y(N760) );
  INVX2TF U577 ( .A(N189), .Y(N780) );
  OAI211X1TF U578 ( .A0(N148), .A1(N777), .B0(N757), .C0(N756), .Y(N758) );
  AOI22X1TF U579 ( .A0(DIVISION_REMA[6]), .A1(N735), .B0(SUM_AB[7]), .B1(N145), 
        .Y(N756) );
  OAI211X1TF U580 ( .A0(N810), .A1(N993), .B0(N755), .C0(N754), .Y(N759) );
  AOI22X1TF U581 ( .A0(X_IN[1]), .A1(N807), .B0(X_IN[0]), .B1(N140), .Y(N754)
         );
  OAI21X1TF U582 ( .A0(N450), .A1(N449), .B0(N459), .Y(N993) );
  OAI22X1TF U583 ( .A0(N189), .A1(N745), .B0(N761), .B1(N154), .Y(N689) );
  AOI211X1TF U584 ( .A0(SUM_AB[5]), .A1(N146), .B0(N744), .C0(N743), .Y(N745)
         );
  OAI211X1TF U585 ( .A0(N810), .A1(N987), .B0(N757), .C0(N742), .Y(N743) );
  OAI21X1TF U586 ( .A0(N429), .A1(N428), .B0(N440), .Y(N987) );
  INVX2TF U587 ( .A(N804), .Y(N791) );
  OAI22X1TF U588 ( .A0(N189), .A1(N734), .B0(N761), .B1(N736), .Y(N691) );
  AOI211X1TF U589 ( .A0(SUM_AB[3]), .A1(N146), .B0(N733), .C0(N732), .Y(N734)
         );
  OAI211X1TF U590 ( .A0(N810), .A1(N981), .B0(N757), .C0(N731), .Y(N732) );
  AOI222X4TF U591 ( .A0(N767), .A1(N105), .B0(N765), .B1(N139), .C0(N557), 
        .C1(N807), .Y(N757) );
  OAI21X1TF U592 ( .A0(N411), .A1(N410), .B0(N419), .Y(N981) );
  OAI22X1TF U593 ( .A0(N730), .A1(N804), .B0(N164), .B1(N104), .Y(N733) );
  NOR3X1TF U594 ( .A(N774), .B(N134), .C(N556), .Y(N782) );
  AOI32X1TF U595 ( .A0(N790), .A1(N816), .A2(N789), .B0(N814), .B1(N156), .Y(
        N685) );
  OAI211X1TF U596 ( .A0(N810), .A1(N999), .B0(N786), .C0(N785), .Y(N787) );
  AOI22X1TF U597 ( .A0(DIVISION_HEAD[1]), .A1(N131), .B0(X_IN[1]), .B1(N105), 
        .Y(N785) );
  OAI21X1TF U598 ( .A0(N475), .A1(N474), .B0(N484), .Y(N999) );
  OAI21X1TF U599 ( .A0(N784), .A1(N804), .B0(N783), .Y(N788) );
  AOI22X1TF U600 ( .A0(DIVISION_REMA[8]), .A1(N134), .B0(N800), .B1(SUM_AB[0]), 
        .Y(N783) );
  AOI22X1TF U601 ( .A0(DIVISION_HEAD[0]), .A1(N806), .B0(SUM_AB[9]), .B1(N146), 
        .Y(N790) );
  OAI22X1TF U602 ( .A0(N510), .A1(N354), .B0(N353), .B1(N352), .Y(N723) );
  AOI211X1TF U603 ( .A0(N491), .A1(N1009), .B0(N350), .C0(N349), .Y(N354) );
  OAI31X1TF U604 ( .A0(XTEMP[12]), .A1(N351), .A2(N506), .B0(N348), .Y(N349)
         );
  INVX2TF U605 ( .A(N608), .Y(N441) );
  NAND2X2TF U606 ( .A(MODE_TYPE[1]), .B(N347), .Y(N608) );
  INVX2TF U607 ( .A(INTADD_0_N1), .Y(N462) );
  NOR2X1TF U608 ( .A(N163), .B(N750), .Y(INTADD_0_CI) );
  INVX2TF U609 ( .A(X_IN[0]), .Y(N750) );
  OAI22X1TF U610 ( .A0(N127), .A1(N1014), .B0(N499), .B1(N102), .Y(N350) );
  NOR2X2TF U611 ( .A(N390), .B(N1014), .Y(N491) );
  AOI31X1TF U612 ( .A0(N84), .A1(N108), .A2(N563), .B0(N344), .Y(N381) );
  OAI211X1TF U613 ( .A0(N108), .A1(N371), .B0(N355), .C0(N343), .Y(N344) );
  NOR2X1TF U614 ( .A(PRE_WORK), .B(N360), .Y(N602) );
  NOR2X1TF U615 ( .A(N367), .B(N944), .Y(N355) );
  INVX2TF U616 ( .A(N390), .Y(N367) );
  INVX2TF U617 ( .A(N617), .Y(N371) );
  AOI32X1TF U618 ( .A0(N817), .A1(N816), .A2(N815), .B0(N814), .B1(N813), .Y(
        N683) );
  AOI211X1TF U619 ( .A0(DIVISION_HEAD[3]), .A1(N131), .B0(N812), .C0(N811), 
        .Y(N815) );
  OAI211X1TF U620 ( .A0(N810), .A1(N1005), .B0(N809), .C0(N808), .Y(N811) );
  AOI22X1TF U621 ( .A0(X_IN[3]), .A1(N105), .B0(X_IN[5]), .B1(N807), .Y(N808)
         );
  AOI22X1TF U622 ( .A0(DIVISION_HEAD[1]), .A1(N134), .B0(DIVISION_HEAD[2]), 
        .B1(N806), .Y(N809) );
  OAI21X1TF U623 ( .A0(N497), .A1(N496), .B0(N1010), .Y(N1005) );
  INVX2TF U624 ( .A(N797), .Y(N810) );
  OAI21X1TF U625 ( .A0(N805), .A1(N804), .B0(N803), .Y(N812) );
  INVX2TF U626 ( .A(N101), .Y(N802) );
  INVX2TF U627 ( .A(N814), .Y(N816) );
  AOI22X1TF U628 ( .A0(N800), .A1(SUM_AB[2]), .B0(SUM_AB[11]), .B1(N146), .Y(
        N817) );
  OAI21X1TF U629 ( .A0(N814), .A1(N555), .B0(N554), .Y(N706) );
  OAI21X1TF U630 ( .A0(N814), .A1(N806), .B0(DIVISION_HEAD[3]), .Y(N554) );
  INVX2TF U631 ( .A(N451), .Y(N806) );
  AOI211X1TF U632 ( .A0(DIVISION_HEAD[2]), .A1(N134), .B0(N553), .C0(N552), 
        .Y(N555) );
  AOI22X1TF U633 ( .A0(N800), .A1(SUM_AB[3]), .B0(N1009), .B1(N797), .Y(N549)
         );
  NOR2X2TF U634 ( .A(N1014), .B(N650), .Y(N797) );
  NOR2X1TF U635 ( .A(N1014), .B(N1010), .Y(N1009) );
  INVX2TF U636 ( .A(SUM_AB[11]), .Y(N496) );
  INVX2TF U637 ( .A(SUM_AB[9]), .Y(N474) );
  INVX2TF U638 ( .A(SUM_AB[7]), .Y(N449) );
  NOR2X1TF U639 ( .A(SUM_AB[6]), .B(N440), .Y(N450) );
  INVX2TF U640 ( .A(SUM_AB[5]), .Y(N428) );
  NOR2X1TF U641 ( .A(SUM_AB[4]), .B(N419), .Y(N429) );
  INVX2TF U642 ( .A(SUM_AB[3]), .Y(N410) );
  NOR3X1TF U643 ( .A(SUM_AB[0]), .B(SUM_AB[2]), .C(SUM_AB[1]), .Y(N411) );
  INVX2TF U644 ( .A(SUM_AB[12]), .Y(N1014) );
  INVX2TF U645 ( .A(N558), .Y(N800) );
  AOI22X1TF U646 ( .A0(N84), .A1(SUM_AB[12]), .B0(X_IN[5]), .B1(N140), .Y(N550) );
  OAI21X1TF U647 ( .A0(N352), .A1(N115), .B0(N253), .Y(OPER_A[12]) );
  AOI22X1TF U648 ( .A0(X_IN[4]), .A1(N106), .B0(X_IN[6]), .B1(N807), .Y(N551)
         );
  AND2X2TF U649 ( .A(N764), .B(N769), .Y(N766) );
  INVX2TF U650 ( .A(N382), .Y(N774) );
  OAI22X1TF U651 ( .A0(N548), .A1(N804), .B0(N547), .B1(N102), .Y(N553) );
  NAND2X2TF U652 ( .A(N347), .B(N307), .Y(N804) );
  AOI32X1TF U653 ( .A0(N84), .A1(N109), .A2(N563), .B0(N617), .B1(N108), .Y(
        N544) );
  INVX2TF U654 ( .A(N347), .Y(N639) );
  AOI31X1TF U655 ( .A0(N122), .A1(N380), .A2(N379), .B0(N378), .Y(N546) );
  INVX2TF U656 ( .A(N302), .Y(N765) );
  OAI211X1TF U657 ( .A0(X_IN[12]), .A1(N547), .B0(N301), .C0(N300), .Y(N302)
         );
  OAI22X1TF U658 ( .A0(Y_IN[10]), .A1(N299), .B0(N298), .B1(N297), .Y(N300) );
  OAI22X1TF U659 ( .A0(X_IN[10]), .A1(N296), .B0(X_IN[11]), .B1(N784), .Y(N297) );
  OAI21X1TF U660 ( .A0(Y_IN[9]), .A1(N295), .B0(Y_IN[8]), .Y(N296) );
  AOI211X1TF U661 ( .A0(X_IN[10]), .A1(N762), .B0(N294), .C0(N293), .Y(N298)
         );
  AOI21X1TF U662 ( .A0(Y_IN[7]), .A1(N498), .B0(N292), .Y(N293) );
  AOI211X1TF U663 ( .A0(X_IN[8]), .A1(N291), .B0(N290), .C0(N289), .Y(N292) );
  NOR2X1TF U664 ( .A(Y_IN[7]), .B(N498), .Y(N290) );
  AOI21X1TF U665 ( .A0(N190), .A1(N466), .B0(N288), .Y(N291) );
  AOI211X1TF U666 ( .A0(X_IN[6]), .A1(N287), .B0(N286), .C0(N285), .Y(N288) );
  NOR2X1TF U667 ( .A(N190), .B(N466), .Y(N286) );
  AOI32X1TF U668 ( .A0(N284), .A1(N283), .A2(N310), .B0(N282), .B1(N283), .Y(
        N287) );
  OAI22X1TF U669 ( .A0(X_IN[4]), .A1(N738), .B0(N107), .B1(N730), .Y(N282) );
  OAI32X1TF U670 ( .A0(N281), .A1(N98), .A2(N308), .B0(X_IN[2]), .B1(N281), 
        .Y(N284) );
  INVX2TF U671 ( .A(X_IN[7]), .Y(N466) );
  INVX2TF U672 ( .A(X_IN[9]), .Y(N498) );
  NOR2X1TF U673 ( .A(Y_IN[9]), .B(N295), .Y(N294) );
  INVX2TF U674 ( .A(X_IN[11]), .Y(N295) );
  NOR2X1TF U675 ( .A(Y_IN[12]), .B(Y_IN[11]), .Y(N301) );
  INVX2TF U676 ( .A(N770), .Y(N557) );
  OR2X2TF U677 ( .A(MODE_TYPE[0]), .B(N307), .Y(N769) );
  INVX2TF U678 ( .A(MODE_TYPE[1]), .Y(N307) );
  OAI31X1TF U679 ( .A0(N277), .A1(N276), .A2(N275), .B0(N274), .Y(N278) );
  NOR2X1TF U680 ( .A(X_IN[10]), .B(N784), .Y(N275) );
  AOI211X1TF U681 ( .A0(X_IN[10]), .A1(N784), .B0(X_IN[9]), .C0(N762), .Y(N276) );
  AOI211X1TF U682 ( .A0(X_IN[9]), .A1(N762), .B0(N273), .C0(N272), .Y(N277) );
  AOI21X1TF U683 ( .A0(Y_IN[7]), .A1(N486), .B0(N271), .Y(N272) );
  AOI211X1TF U684 ( .A0(N270), .A1(X_IN[7]), .B0(N269), .C0(N268), .Y(N271) );
  NOR2X1TF U685 ( .A(Y_IN[7]), .B(N486), .Y(N269) );
  AOI21X1TF U686 ( .A0(N190), .A1(N460), .B0(N267), .Y(N270) );
  AOI211X1TF U687 ( .A0(N266), .A1(X_IN[5]), .B0(N265), .C0(N264), .Y(N267) );
  NOR2X1TF U688 ( .A(N190), .B(N460), .Y(N265) );
  AOI211X1TF U689 ( .A0(Y_IN[3]), .A1(N438), .B0(N263), .C0(N262), .Y(N266) );
  AOI211X1TF U690 ( .A0(X_IN[4]), .A1(N730), .B0(N98), .C0(N738), .Y(N262) );
  OAI32X1TF U691 ( .A0(N261), .A1(X_IN[2]), .A2(N308), .B0(X_IN[1]), .B1(N261), 
        .Y(N263) );
  OAI211X1TF U692 ( .A0(Y_IN[3]), .A1(N438), .B0(N260), .C0(N310), .Y(N261) );
  AOI22X1TF U693 ( .A0(N98), .A1(N738), .B0(X_IN[2]), .B1(N309), .Y(N260) );
  INVX2TF U694 ( .A(X_IN[4]), .Y(N438) );
  INVX2TF U695 ( .A(X_IN[6]), .Y(N460) );
  INVX2TF U696 ( .A(X_IN[8]), .Y(N486) );
  NOR2X1TF U697 ( .A(Y_IN[9]), .B(N499), .Y(N273) );
  INVX2TF U698 ( .A(X_IN[10]), .Y(N499) );
  NOR2X1TF U699 ( .A(Y_IN[11]), .B(N299), .Y(N279) );
  INVX2TF U700 ( .A(X_IN[12]), .Y(N299) );
  INVX2TF U701 ( .A(N333), .Y(N380) );
  OAI211X1TF U702 ( .A0(N849), .A1(N848), .B0(N847), .C0(N846), .Y(N678) );
  AOI32X1TF U703 ( .A0(N932), .A1(OPER_B[4]), .A2(N845), .B0(N877), .B1(
        OPER_B[4]), .Y(N846) );
  AOI211X1TF U704 ( .A0(N851), .A1(OPER_B[5]), .B0(N844), .C0(N843), .Y(N847)
         );
  OAI31X1TF U705 ( .A0(N929), .A1(OPER_A[4]), .A2(N842), .B0(N201), .Y(N843)
         );
  AOI21X1TF U706 ( .A0(N116), .A1(C152_DATA4_4), .B0(N202), .Y(N201) );
  NOR3X1TF U707 ( .A(OPER_B[4]), .B(N845), .C(N119), .Y(N844) );
  AOI21X1TF U708 ( .A0(N926), .A1(N842), .B0(N841), .Y(N848) );
  INVX2TF U709 ( .A(N927), .Y(N841) );
  AOI211X1TF U710 ( .A0(N117), .A1(C152_DATA4_5), .B0(N853), .C0(N207), .Y(
        N208) );
  OAI31X1TF U711 ( .A0(OPER_B[5]), .A1(N852), .A2(N119), .B0(N892), .Y(N853)
         );
  OAI211X1TF U712 ( .A0(SIGN_Y), .A1(N961), .B0(N217), .C0(N968), .Y(N892) );
  AOI22X1TF U713 ( .A0(N851), .A1(OPER_B[6]), .B0(N850), .B1(N855), .Y(N860)
         );
  NOR2X1TF U714 ( .A(N929), .B(OPER_A[5]), .Y(N850) );
  INVX2TF U715 ( .A(N881), .Y(N851) );
  AOI22X1TF U716 ( .A0(OPER_B[5]), .A1(N857), .B0(OPER_A[5]), .B1(N856), .Y(
        N859) );
  OAI21X1TF U717 ( .A0(N929), .A1(N855), .B0(N927), .Y(N856) );
  OAI21X1TF U718 ( .A0(N119), .A1(N854), .B0(N930), .Y(N857) );
  AOI22X1TF U719 ( .A0(OPER_B[9]), .A1(N900), .B0(OPER_A[9]), .B1(N899), .Y(
        N901) );
  OAI21X1TF U720 ( .A0(N929), .A1(N898), .B0(N927), .Y(N899) );
  OAI21X1TF U721 ( .A0(N119), .A1(N897), .B0(N930), .Y(N900) );
  AOI31X1TF U722 ( .A0(N932), .A1(N186), .A2(N897), .B0(N896), .Y(N902) );
  OAI211X1TF U723 ( .A0(N170), .A1(N939), .B0(N204), .C0(N203), .Y(N896) );
  AOI22X1TF U724 ( .A0(SIGN_Y), .A1(N894), .B0(N893), .B1(N898), .Y(N903) );
  NOR2X1TF U725 ( .A(N929), .B(OPER_A[9]), .Y(N893) );
  OR2X2TF U726 ( .A(N924), .B(N878), .Y(N202) );
  NOR2X1TF U727 ( .A(N963), .B(N829), .Y(N863) );
  INVX2TF U728 ( .A(N930), .Y(N877) );
  OAI211X1TF U729 ( .A0(N185), .A1(N939), .B0(N938), .C0(N937), .Y(N671) );
  AOI211X1TF U730 ( .A0(OPER_A[11]), .A1(N936), .B0(N935), .C0(N934), .Y(N937)
         );
  AOI21X1TF U731 ( .A0(N960), .A1(N217), .B0(N205), .Y(N206) );
  NOR3X1TF U732 ( .A(N118), .B(OPER_B[11]), .C(N933), .Y(N205) );
  INVX2TF U733 ( .A(N931), .Y(N933) );
  NOR3X1TF U734 ( .A(N108), .B(N176), .C(N961), .Y(N960) );
  OAI22X1TF U735 ( .A0(N136), .A1(N198), .B0(N125), .B1(OFFSET[2]), .Y(C2_Z_4)
         );
  INVX2TF U736 ( .A(Y_IN[4]), .Y(N198) );
  OAI22X1TF U737 ( .A0(N136), .A1(N197), .B0(N125), .B1(OFFSET[3]), .Y(C2_Z_5)
         );
  OAI22X1TF U738 ( .A0(N136), .A1(N196), .B0(N125), .B1(OFFSET[4]), .Y(C2_Z_6)
         );
  OAI22X1TF U739 ( .A0(N135), .A1(N191), .B0(N125), .B1(OFFSET[5]), .Y(C2_Z_7)
         );
  OAI22X1TF U740 ( .A0(N136), .A1(N762), .B0(N125), .B1(OFFSET[6]), .Y(C2_Z_8)
         );
  OAI22X1TF U741 ( .A0(N135), .A1(N784), .B0(N125), .B1(OFFSET[7]), .Y(C2_Z_9)
         );
  OAI22X1TF U742 ( .A0(N136), .A1(N547), .B0(N125), .B1(OFFSET[8]), .Y(C2_Z_10) );
  OAI22X1TF U743 ( .A0(N136), .A1(N805), .B0(N125), .B1(OFFSET[9]), .Y(C2_Z_11) );
  INVX2TF U744 ( .A(Y_IN[11]), .Y(N805) );
  OAI32X1TF U745 ( .A0(N183), .A1(N931), .A2(N119), .B0(N930), .B1(N183), .Y(
        N935) );
  NOR2X1TF U746 ( .A(OPER_B[9]), .B(N897), .Y(N917) );
  NOR2X1TF U747 ( .A(N862), .B(OPER_B[6]), .Y(N879) );
  INVX2TF U748 ( .A(N866), .Y(N862) );
  NOR2X1TF U749 ( .A(OPER_B[5]), .B(N854), .Y(N866) );
  NOR2X1TF U750 ( .A(OPER_B[3]), .B(N834), .Y(N845) );
  OAI21X1TF U751 ( .A0(N929), .A1(N928), .B0(N927), .Y(N936) );
  AOI31X1TF U752 ( .A0(N926), .A1(N925), .A2(N928), .B0(N924), .Y(N938) );
  AOI211X1TF U753 ( .A0(N109), .A1(N961), .B0(SIGN_Y), .C0(N904), .Y(N924) );
  NOR2X1TF U754 ( .A(OPER_A[9]), .B(N898), .Y(N911) );
  NOR2X1TF U755 ( .A(OPER_A[7]), .B(N880), .Y(N885) );
  NOR2X1TF U756 ( .A(OPER_A[5]), .B(N855), .Y(N869) );
  NOR2X1TF U757 ( .A(OPER_A[3]), .B(N833), .Y(N842) );
  OAI21X1TF U758 ( .A0(N520), .A1(N115), .B0(N244), .Y(OPER_A[4]) );
  OAI21X1TF U759 ( .A0(N439), .A1(N115), .B0(N245), .Y(OPER_A[5]) );
  OAI21X1TF U760 ( .A0(N525), .A1(N115), .B0(N246), .Y(OPER_A[6]) );
  OAI21X1TF U761 ( .A0(N461), .A1(N115), .B0(N247), .Y(OPER_A[7]) );
  OAI21X1TF U762 ( .A0(N159), .A1(N115), .B0(N248), .Y(OPER_A[8]) );
  OAI21X1TF U763 ( .A0(N115), .A1(N528), .B0(N249), .Y(OPER_A[9]) );
  OAI21X1TF U764 ( .A0(N115), .A1(N160), .B0(N250), .Y(OPER_A[10]) );
  OAI21X1TF U765 ( .A0(N115), .A1(N153), .B0(N251), .Y(OPER_A[11]) );
  OAI211X1TF U766 ( .A0(N175), .A1(N939), .B0(N840), .C0(N839), .Y(N679) );
  AOI211X1TF U767 ( .A0(OPER_A[3]), .A1(N838), .B0(N837), .C0(N836), .Y(N839)
         );
  OAI31X1TF U768 ( .A0(N929), .A1(OPER_A[3]), .A2(N835), .B0(N200), .Y(N836)
         );
  AOI21X1TF U769 ( .A0(C152_DATA4_3), .A1(N116), .B0(N894), .Y(N200) );
  OAI21X1TF U770 ( .A0(N136), .A1(N308), .B0(N120), .Y(C2_Z_1) );
  OAI22X1TF U771 ( .A0(N136), .A1(N730), .B0(N120), .B1(OFFSET[1]), .Y(C2_Z_3)
         );
  INVX2TF U772 ( .A(Y_IN[3]), .Y(N730) );
  OAI32X1TF U773 ( .A0(N181), .A1(N118), .A2(N834), .B0(N930), .B1(N181), .Y(
        N837) );
  INVX2TF U774 ( .A(N861), .Y(N915) );
  AOI32X1TF U775 ( .A0(N605), .A1(N341), .A2(N824), .B0(N946), .B1(N340), .Y(
        N861) );
  INVX2TF U776 ( .A(N941), .Y(N946) );
  OAI21X1TF U777 ( .A0(N929), .A1(N833), .B0(N927), .Y(N838) );
  INVX2TF U778 ( .A(N830), .Y(N906) );
  AOI21X1TF U779 ( .A0(N564), .A1(N340), .B0(N563), .Y(N830) );
  INVX2TF U780 ( .A(N835), .Y(N833) );
  NOR3X1TF U781 ( .A(OPER_A[2]), .B(OPER_A[1]), .C(OPER_A[0]), .Y(N835) );
  OAI21X1TF U782 ( .A0(N151), .A1(N114), .B0(N242), .Y(OPER_A[2]) );
  INVX2TF U783 ( .A(N926), .Y(N929) );
  NOR2X2TF U784 ( .A(N918), .B(N910), .Y(N926) );
  INVX2TF U785 ( .A(N891), .Y(N918) );
  OAI21X1TF U786 ( .A0(N152), .A1(N114), .B0(N243), .Y(OPER_A[3]) );
  AOI31X1TF U787 ( .A0(N932), .A1(N181), .A2(N834), .B0(N875), .Y(N840) );
  OAI21X1TF U788 ( .A0(N971), .A1(N904), .B0(N832), .Y(N875) );
  INVX2TF U789 ( .A(N904), .Y(N217) );
  INVX2TF U790 ( .A(N339), .Y(N955) );
  INVX2TF U791 ( .A(N565), .Y(N948) );
  NOR2X1TF U792 ( .A(OPER_B[1]), .B(OPER_B[0]), .Y(N831) );
  AOI22X1TF U793 ( .A0(N108), .A1(DIVISION_HEAD[3]), .B0(XTEMP[12]), .B1(N109), 
        .Y(N340) );
  INVX2TF U794 ( .A(N605), .Y(N823) );
  NOR2X2TF U795 ( .A(N603), .B(N631), .Y(N824) );
  AOI221X1TF U796 ( .A0(N128), .A1(N167), .B0(N179), .B1(N91), .C0(N819), .Y(
        N820) );
  AOI22X1TF U797 ( .A0(\INDEX[2] ), .A1(N90), .B0(N124), .B1(\RSHT_BITS[3] ), 
        .Y(N818) );
  AOI32X1TF U798 ( .A0(N941), .A1(N949), .A2(N364), .B0(N951), .B1(N949), .Y(
        N337) );
  OR2X2TF U799 ( .A(N631), .B(N161), .Y(N364) );
  INVX2TF U800 ( .A(N603), .Y(N642) );
  OAI21X1TF U801 ( .A0(N339), .A1(N940), .B0(N335), .Y(N607) );
  OAI21X1TF U802 ( .A0(N570), .A1(N564), .B0(N336), .Y(N335) );
  NOR2X2TF U803 ( .A(\RSHT_BITS[3] ), .B(N591), .Y(N605) );
  NOR3X1TF U804 ( .A(N121), .B(N122), .C(N950), .Y(N822) );
  NOR2X1TF U805 ( .A(SIGN_Y), .B(N63), .Y(N895) );
  INVX2TF U806 ( .A(N306), .Y(N627) );
  OAI22X1TF U807 ( .A0(Y_IN[12]), .A1(N159), .B0(N331), .B1(N330), .Y(N332) );
  OAI31X1TF U808 ( .A0(N329), .A1(DIVISION_HEAD[10]), .A2(N547), .B0(N328), 
        .Y(N330) );
  AOI22X1TF U809 ( .A0(Y_IN[11]), .A1(N461), .B0(N327), .B1(N326), .Y(N328) );
  OAI22X1TF U810 ( .A0(DIVISION_HEAD[8]), .A1(N762), .B0(DIVISION_HEAD[9]), 
        .B1(N784), .Y(N326) );
  INVX2TF U811 ( .A(N325), .Y(N327) );
  NOR2X1TF U812 ( .A(Y_IN[11]), .B(N461), .Y(N329) );
  AOI211X1TF U813 ( .A0(DIVISION_HEAD[8]), .A1(N762), .B0(N324), .C0(N325), 
        .Y(N331) );
  OAI21X1TF U814 ( .A0(Y_IN[11]), .A1(N461), .B0(N323), .Y(N325) );
  INVX2TF U815 ( .A(Y_IN[9]), .Y(N784) );
  INVX2TF U816 ( .A(Y_IN[10]), .Y(N547) );
  AOI21X1TF U817 ( .A0(N97), .A1(N152), .B0(N322), .Y(N324) );
  AOI211X1TF U818 ( .A0(N321), .A1(DIVISION_HEAD[6]), .B0(N320), .C0(N319), 
        .Y(N322) );
  NOR2X1TF U819 ( .A(N97), .B(N152), .Y(N320) );
  AOI211X1TF U820 ( .A0(N317), .A1(DIVISION_HEAD[4]), .B0(N316), .C0(N315), 
        .Y(N318) );
  NOR2X1TF U821 ( .A(Y_IN[5]), .B(N511), .Y(N316) );
  AOI21X1TF U822 ( .A0(Y_IN[3]), .A1(N648), .B0(N314), .Y(N317) );
  OAI32X1TF U823 ( .A0(N313), .A1(DIVISION_HEAD[2]), .A2(N738), .B0(N312), 
        .B1(N313), .Y(N314) );
  OAI211X1TF U824 ( .A0(Y_IN[2]), .A1(N813), .B0(N311), .C0(N310), .Y(N312) );
  INVX2TF U825 ( .A(Y_IN[0]), .Y(N656) );
  INVX2TF U826 ( .A(Y_IN[1]), .Y(N308) );
  INVX2TF U827 ( .A(Y_IN[2]), .Y(N738) );
  INVX2TF U828 ( .A(Y_IN[8]), .Y(N762) );
  INVX2TF U829 ( .A(Y_IN[12]), .Y(N548) );
  NOR2X1TF U830 ( .A(N238), .B(N352), .Y(FOUT[12]) );
  AND2X2TF U831 ( .A(ZTEMP[12]), .B(N143), .Y(POUT[12]) );
  OAI21X1TF U832 ( .A0(N151), .A1(N238), .B0(N223), .Y(FOUT[2]) );
  AOI21X1TF U833 ( .A0(N216), .A1(DIVISION_REMA[2]), .B0(N222), .Y(N223) );
  OAI22X1TF U834 ( .A0(N520), .A1(N94), .B0(N157), .B1(N88), .Y(N222) );
  AND2X2TF U835 ( .A(ZTEMP[2]), .B(N188), .Y(POUT[2]) );
  AND2X2TF U836 ( .A(ZTEMP[10]), .B(N143), .Y(POUT[10]) );
  OAI21X1TF U837 ( .A0(N152), .A1(N238), .B0(N225), .Y(FOUT[3]) );
  AOI21X1TF U838 ( .A0(N216), .A1(DIVISION_REMA[3]), .B0(N224), .Y(N225) );
  OAI22X1TF U839 ( .A0(N439), .A1(N93), .B0(N154), .B1(N88), .Y(N224) );
  AND2X2TF U840 ( .A(ZTEMP[3]), .B(N188), .Y(POUT[3]) );
  AND2X2TF U841 ( .A(ZTEMP[9]), .B(N143), .Y(POUT[9]) );
  NOR2X1TF U842 ( .A(N238), .B(N153), .Y(FOUT[11]) );
  AND2X2TF U843 ( .A(ZTEMP[11]), .B(N143), .Y(POUT[11]) );
  OAI21X1TF U844 ( .A0(N159), .A1(N238), .B0(N235), .Y(FOUT[8]) );
  AOI21X1TF U845 ( .A0(N216), .A1(DIVISION_REMA[8]), .B0(N234), .Y(N235) );
  OAI22X1TF U846 ( .A0(N149), .A1(N89), .B0(N160), .B1(N93), .Y(N234) );
  AND2X2TF U847 ( .A(ZTEMP[8]), .B(N143), .Y(POUT[8]) );
  OAI21X1TF U848 ( .A0(N511), .A1(N238), .B0(N221), .Y(FOUT[1]) );
  AOI21X1TF U849 ( .A0(N216), .A1(DIVISION_REMA[1]), .B0(N220), .Y(N221) );
  OAI22X1TF U850 ( .A0(N152), .A1(N93), .B0(N736), .B1(N88), .Y(N220) );
  AND2X2TF U851 ( .A(ZTEMP[1]), .B(N188), .Y(POUT[1]) );
  OAI21X1TF U852 ( .A0(N439), .A1(N238), .B0(N229), .Y(FOUT[5]) );
  AOI21X1TF U853 ( .A0(N216), .A1(DIVISION_REMA[5]), .B0(N228), .Y(N229) );
  OAI22X1TF U854 ( .A0(N461), .A1(N93), .B0(N155), .B1(N88), .Y(N228) );
  OAI21X1TF U855 ( .A0(N520), .A1(N141), .B0(N227), .Y(FOUT[4]) );
  AOI21X1TF U856 ( .A0(N216), .A1(DIVISION_REMA[4]), .B0(N226), .Y(N227) );
  OAI22X1TF U857 ( .A0(N525), .A1(N94), .B0(N158), .B1(N88), .Y(N226) );
  AND2X2TF U858 ( .A(ZTEMP[4]), .B(N188), .Y(POUT[4]) );
  OAI21X1TF U859 ( .A0(N461), .A1(N238), .B0(N233), .Y(FOUT[7]) );
  AOI21X1TF U860 ( .A0(N216), .A1(DIVISION_REMA[7]), .B0(N232), .Y(N233) );
  OAI22X1TF U861 ( .A0(N156), .A1(N89), .B0(N528), .B1(N93), .Y(N232) );
  OAI21X1TF U862 ( .A0(N525), .A1(N141), .B0(N231), .Y(FOUT[6]) );
  AOI21X1TF U863 ( .A0(N216), .A1(DIVISION_REMA[6]), .B0(N230), .Y(N231) );
  OAI22X1TF U864 ( .A0(N159), .A1(N94), .B0(N148), .B1(N89), .Y(N230) );
  INVX2TF U865 ( .A(N256), .Y(N238) );
  NOR2X1TF U866 ( .A(N333), .B(N365), .Y(ALU_IS_DONE) );
  OAI211X1TF U867 ( .A0(N151), .A1(N94), .B0(N219), .C0(N218), .Y(FOUT[0]) );
  AND2X2TF U868 ( .A(ZTEMP[0]), .B(N143), .Y(POUT[0]) );
  AOI22X1TF U869 ( .A0(N133), .A1(\INTADD_0_SUM[5] ), .B0(N800), .B1(
        SUM_AB[10]), .Y(N445) );
  AOI21X1TF U870 ( .A0(N133), .A1(N470), .B0(N469), .Y(N471) );
  AOI22X1TF U871 ( .A0(N132), .A1(N463), .B0(SUM_AB[8]), .B1(N137), .Y(N465)
         );
  AOI22X1TF U872 ( .A0(N133), .A1(\INTADD_0_SUM[3] ), .B0(SUM_AB[4]), .B1(N138), .Y(N427) );
  AOI22X1TF U873 ( .A0(N133), .A1(\INTADD_0_SUM[1] ), .B0(SUM_AB[2]), .B1(N138), .Y(N408) );
  AOI31X1TF U874 ( .A0(X_IN[0]), .A1(N133), .A2(N163), .B0(N386), .Y(N387) );
  AOI22X1TF U875 ( .A0(N133), .A1(\INTADD_0_SUM[0] ), .B0(SUM_AB[1]), .B1(N138), .Y(N398) );
  AOI22X1TF U876 ( .A0(N133), .A1(\INTADD_0_SUM[6] ), .B0(SUM_AB[7]), .B1(N138), .Y(N458) );
  AOI22X1TF U877 ( .A0(N132), .A1(\INTADD_0_SUM[4] ), .B0(SUM_AB[5]), .B1(N137), .Y(N434) );
  AOI31X1TF U878 ( .A0(N132), .A1(N160), .A2(N492), .B0(N487), .Y(N488) );
  AOI22X1TF U879 ( .A0(N133), .A1(\INTADD_0_SUM[2] ), .B0(SUM_AB[3]), .B1(N138), .Y(N418) );
  AOI31X1TF U880 ( .A0(N133), .A1(N153), .A2(N507), .B0(N505), .Y(N509) );
  AOI21X1TF U881 ( .A0(N133), .A1(N351), .B0(N510), .Y(N353) );
  NAND3X1TF U882 ( .A(N892), .B(N211), .C(N210), .Y(N674) );
  OAI2BB1X1TF U883 ( .A0N(N117), .A1N(C152_DATA4_10), .B0(N212), .Y(N672) );
  NAND3X1TF U884 ( .A(N859), .B(N860), .C(N208), .Y(N677) );
  OR3X1TF U885 ( .A(N904), .B(N74), .C(N895), .Y(N203) );
  NAND2X1TF U886 ( .A(N116), .B(C152_DATA4_9), .Y(N204) );
  OAI2BB1X1TF U887 ( .A0N(N116), .A1N(C152_DATA4_11), .B0(N206), .Y(N934) );
  NAND2BX1TF U888 ( .AN(DP_OP_333_124_4748_N57), .B(N135), .Y(N199) );
  OAI2BB2XLTF U889 ( .B0(OFFSET[0]), .B1(N120), .A0N(Y_IN[2]), .A1N(N967), .Y(
        C2_Z_2) );
  INVX2TF U890 ( .A(N956), .Y(N963) );
  AOI2BB2X1TF U891 ( .B0(N216), .B1(DIVISION_REMA[0]), .A0N(N164), .A1N(N89), 
        .Y(N219) );
  OAI222X1TF U892 ( .A0(N94), .A1(N352), .B0(N89), .B1(N648), .C0(N238), .C1(
        N160), .Y(FOUT[10]) );
  OAI222X1TF U893 ( .A0(N238), .A1(N528), .B0(N89), .B1(N813), .C0(N153), .C1(
        N94), .Y(FOUT[9]) );
  NAND2X1TF U894 ( .A(N161), .B(N172), .Y(N365) );
  NAND3X1TF U895 ( .A(STEP[2]), .B(STEP[3]), .C(N642), .Y(N941) );
  NAND3X1TF U896 ( .A(N545), .B(N382), .C(N634), .Y(N647) );
  NOR4XLTF U897 ( .A(N763), .B(N617), .C(N802), .D(N647), .Y(N259) );
  AOI222XLTF U898 ( .A0(STEP[2]), .A1(N162), .B0(N121), .B1(N172), .C0(N150), 
        .C1(N122), .Y(N257) );
  NAND3X1TF U899 ( .A(N259), .B(N356), .C(N633), .Y(N619) );
  NAND2X1TF U900 ( .A(Y_IN[1]), .B(Y_IN[0]), .Y(N309) );
  AOI2BB1X1TF U901 ( .A0N(X_IN[5]), .A1N(N266), .B0(Y_IN[4]), .Y(N264) );
  AOI2BB1X1TF U902 ( .A0N(X_IN[7]), .A1N(N270), .B0(Y_IN[6]), .Y(N268) );
  NAND2X1TF U903 ( .A(MODE_TYPE[0]), .B(N307), .Y(N764) );
  AO22X1TF U904 ( .A0(X_IN[4]), .A1(N738), .B0(N98), .B1(N309), .Y(N281) );
  NAND2X1TF U905 ( .A(N107), .B(N730), .Y(N283) );
  AOI2BB1X1TF U906 ( .A0N(N287), .A1N(X_IN[6]), .B0(Y_IN[4]), .Y(N285) );
  AOI2BB1X1TF U907 ( .A0N(N291), .A1N(X_IN[8]), .B0(Y_IN[6]), .Y(N289) );
  NAND2X1TF U908 ( .A(N166), .B(N179), .Y(N616) );
  NAND2X1TF U909 ( .A(N831), .B(N165), .Y(N834) );
  NAND2X1TF U910 ( .A(N845), .B(N175), .Y(N854) );
  NOR2BX1TF U911 ( .AN(N879), .B(OPER_B[7]), .Y(N882) );
  NAND2X1TF U912 ( .A(N882), .B(N169), .Y(N897) );
  NAND2X1TF U913 ( .A(N917), .B(N170), .Y(N931) );
  NAND2X1TF U914 ( .A(N895), .B(N74), .Y(N954) );
  NAND2X1TF U915 ( .A(N565), .B(N954), .Y(N940) );
  NAND2X1TF U916 ( .A(N963), .B(N373), .Y(N573) );
  NAND3X1TF U917 ( .A(N92), .B(N91), .C(N90), .Y(N591) );
  NOR2BX1TF U918 ( .AN(N573), .B(N605), .Y(N570) );
  NAND2X1TF U919 ( .A(PRE_WORK), .B(N345), .Y(N949) );
  NAND2X1TF U920 ( .A(N605), .B(N824), .Y(N338) );
  NAND2X1TF U921 ( .A(N215), .B(N955), .Y(N358) );
  NAND3X1TF U922 ( .A(SIGN_Y), .B(N74), .C(N894), .Y(N825) );
  NAND2X1TF U923 ( .A(N849), .B(N842), .Y(N855) );
  NAND2X1TF U924 ( .A(N868), .B(N869), .Y(N880) );
  NAND2X1TF U925 ( .A(N884), .B(N885), .Y(N898) );
  NAND2X1TF U926 ( .A(N909), .B(N911), .Y(N928) );
  NAND3X1TF U927 ( .A(N605), .B(N602), .C(N171), .Y(N600) );
  NAND2X1TF U928 ( .A(N411), .B(N410), .Y(N419) );
  NAND2X1TF U929 ( .A(N429), .B(N428), .Y(N440) );
  NAND2X1TF U930 ( .A(N450), .B(N449), .Y(N459) );
  NAND2X1TF U931 ( .A(N497), .B(N496), .Y(N1010) );
  AOI222XLTF U932 ( .A0(XTEMP[11]), .A1(X_IN[11]), .B0(XTEMP[11]), .B1(N495), 
        .C0(X_IN[11]), .C1(N495), .Y(N346) );
  XOR2X1TF U933 ( .A(X_IN[12]), .B(N346), .Y(N351) );
  NAND3X1TF U934 ( .A(N566), .B(POST_WORK), .C(N602), .Y(N368) );
  NAND3BX1TF U935 ( .AN(N358), .B(N948), .C(N963), .Y(N598) );
  NAND3X1TF U936 ( .A(N609), .B(N359), .C(N598), .Y(N943) );
  NAND2X1TF U937 ( .A(N127), .B(N390), .Y(N377) );
  NAND3X1TF U938 ( .A(N380), .B(N122), .C(DP_OP_333_124_4748_N57), .Y(N638) );
  NOR2BX1TF U939 ( .AN(N634), .B(N944), .Y(N542) );
  NAND3X1TF U940 ( .A(N542), .B(N372), .C(N371), .Y(N376) );
  NAND4X1TF U941 ( .A(N423), .B(N422), .C(N421), .D(N420), .Y(N424) );
  NAND4X1TF U942 ( .A(N434), .B(N433), .C(N432), .D(N431), .Y(N435) );
  NAND4X1TF U943 ( .A(N445), .B(N444), .C(N443), .D(N442), .Y(N446) );
  OAI2BB1X1TF U944 ( .A0N(DIVISION_HEAD[10]), .A1N(N469), .B0(N448), .Y(N713)
         );
  AOI2BB2X1TF U945 ( .B0(X_IN[9]), .B1(N476), .A0N(N476), .A1N(X_IN[9]), .Y(
        N481) );
  NAND3X1TF U946 ( .A(N132), .B(N528), .C(N481), .Y(N477) );
  AOI2BB1X1TF U947 ( .A0N(N506), .A1N(N481), .B0(N510), .Y(N482) );
  AOI2BB2X1TF U948 ( .B0(N485), .B1(N499), .A0N(N499), .A1N(N485), .Y(N492) );
  AOI2BB1X1TF U949 ( .A0N(N506), .A1N(N492), .B0(N510), .Y(N493) );
  AOI2BB2X1TF U950 ( .B0(N86), .B1(N495), .A0N(N495), .A1N(N86), .Y(N507) );
  OAI2BB2XLTF U951 ( .B0(N499), .B1(N608), .A0N(XTEMP[12]), .A1N(N99), .Y(N500) );
  AOI2BB1X1TF U952 ( .A0N(N506), .A1N(N507), .B0(N510), .Y(N508) );
  AOI2BB1X1TF U953 ( .A0N(DIVISION_REMA[2]), .A1N(N515), .B0(DIVISION_HEAD[6]), 
        .Y(N513) );
  OA21XLTF U954 ( .A0(N520), .A1(DIVISION_REMA[4]), .B0(N517), .Y(N519) );
  OA21XLTF U955 ( .A0(N525), .A1(DIVISION_REMA[6]), .B0(N522), .Y(N524) );
  OA21XLTF U956 ( .A0(XTEMP[12]), .A1(N535), .B0(N648), .Y(N534) );
  NAND4X1TF U957 ( .A(N545), .B(N544), .C(N638), .D(N543), .Y(N556) );
  NAND3X1TF U958 ( .A(N551), .B(N550), .C(N549), .Y(N552) );
  NAND3X1TF U959 ( .A(N757), .B(N559), .C(N558), .Y(N560) );
  NAND3X1TF U960 ( .A(N566), .B(N602), .C(N823), .Y(N572) );
  NAND4X1TF U961 ( .A(N568), .B(N567), .C(N639), .D(N572), .Y(N569) );
  NAND2X1TF U962 ( .A(N178), .B(N167), .Y(N590) );
  NOR4XLTF U963 ( .A(\RSHT_BITS[3] ), .B(N90), .C(N614), .D(N590), .Y(N571) );
  NAND2X1TF U964 ( .A(N579), .B(N589), .Y(N586) );
  NAND2X1TF U965 ( .A(N92), .B(N91), .Y(N588) );
  AOI2BB2X1TF U966 ( .B0(N596), .B1(N167), .A0N(N590), .A1N(N592), .Y(N584) );
  NAND4X1TF U967 ( .A(N104), .B(N634), .C(N633), .D(N632), .Y(N635) );
  NAND4X1TF U968 ( .A(N640), .B(N639), .C(N638), .D(N643), .Y(N697) );
  NAND3X1TF U969 ( .A(N757), .B(N652), .C(N651), .Y(N653) );
  AO22X1TF U970 ( .A0(DIVISION_REMA[4]), .A1(N735), .B0(N190), .B1(N791), .Y(
        N744) );
  AOI2BB1X1TF U971 ( .A0N(X_IN[1]), .A1N(N765), .B0(N764), .Y(N768) );
  NAND4X1TF U972 ( .A(N795), .B(N794), .C(N793), .D(N792), .Y(N796) );
  OAI221XLTF U973 ( .A0(\INDEX[2] ), .A1(N90), .B0(N124), .B1(\RSHT_BITS[3] ), 
        .C0(N818), .Y(N819) );
  OAI221XLTF U974 ( .A0(N129), .A1(N178), .B0(N166), .B1(N92), .C0(N820), .Y(
        N829) );
  NAND2X1TF U975 ( .A(N891), .B(N863), .Y(N858) );
  NAND2BX1TF U976 ( .AN(N821), .B(N858), .Y(N878) );
  NAND2X1TF U977 ( .A(N828), .B(N963), .Y(N864) );
  NAND3X1TF U978 ( .A(SIGN_Y), .B(N74), .C(N217), .Y(N832) );
  OAI2BB1X1TF U979 ( .A0N(N956), .A1N(N829), .B0(N828), .Y(N914) );
  NAND3X1TF U980 ( .A(N74), .B(N176), .C(N109), .Y(N971) );
  NAND2X1TF U981 ( .A(N891), .B(N914), .Y(N939) );
  NAND3X1TF U982 ( .A(N903), .B(N902), .C(N901), .Y(N673) );
  NAND2X1TF U983 ( .A(N975), .B(N974), .Y(N668) );
  NAND2X1TF U984 ( .A(N978), .B(N977), .Y(N667) );
  NAND2X1TF U985 ( .A(SUM_AB[3]), .B(N96), .Y(N979) );
  NAND2X1TF U986 ( .A(N984), .B(N983), .Y(N665) );
  NAND2X1TF U987 ( .A(SUM_AB[5]), .B(N96), .Y(N985) );
  NAND2X1TF U988 ( .A(N990), .B(N989), .Y(N663) );
  NAND2X1TF U989 ( .A(SUM_AB[7]), .B(N96), .Y(N991) );
  NAND2X1TF U990 ( .A(N996), .B(N995), .Y(N661) );
  NAND2X1TF U991 ( .A(SUM_AB[9]), .B(N96), .Y(N997) );
  NAND2X1TF U992 ( .A(N1002), .B(N1001), .Y(N659) );
  NAND2X1TF U993 ( .A(SUM_AB[11]), .B(N96), .Y(N1003) );
endmodule


module SERIAL_CPU_8BIT_VG ( CLK, ENABLE, RST_N, START, I_DATAIN, D_DATAIN, 
        IS_I_ADDR, NXT, I_ADDR, D_ADDR, D_WE, D_DATAOUT, IO_STATUS, IO_CONTROL, 
        IO_DATAINA, IO_DATAINB, IO_DATAOUTA, IO_DATAOUTB, IO_OFFSET );
  input [7:0] I_DATAIN;
  input [7:0] D_DATAIN;
  output [1:0] NXT;
  output [8:0] I_ADDR;
  output [8:0] D_ADDR;
  output [7:0] D_DATAOUT;
  input [15:0] IO_STATUS;
  output [15:0] IO_CONTROL;
  input [15:0] IO_DATAINA;
  input [15:0] IO_DATAINB;
  output [15:0] IO_DATAOUTA;
  output [15:0] IO_DATAOUTB;
  output [15:0] IO_OFFSET;
  input CLK, ENABLE, RST_N, START;
  output IS_I_ADDR, D_WE;
  wire   \OPER1_R1[2] , N114, N162, N163, N164, CF_BUF, N466, N467, N468, N469,
         N470, N471, N472, N473, N474, N475, N476, N477, N478, N479, N480,
         N481, N482, N500, N501, N502, N503, N504, N505, N506, N507, N508,
         N509, N510, N511, N512, N513, N514, N515, N516, N584, N585, ZF, NF,
         CF, N612, N412, N414, N415, N416, N417, N418, N420, N421, N423, N424,
         N429, N431, N432, N442, N443, N444, N445, N446, N447, N448, N449,
         N450, N451, N452, N453, N454, N455, N456, N457, N458, N460, N461,
         N462, N463, N464, N465, N4660, N4670, N4680, N4690, N4700, N4710,
         N4720, N4730, N4740, N4750, N4760, N4770, N4780, N4790, N4800, N4810,
         N4820, N483, N484, N485, N486, N487, N488, N492, N493, N494, N495,
         N496, N497, N498, N499, N5030, N5040, N5060, N5070, N5090, N5100,
         N5120, N5130, N5150, N5160, N518, N519, N521, N522, N524, N525, N527,
         N528, N530, N531, N533, N534, N536, N537, N539, N540, N542, N543,
         N545, N558, N562, N564, N579, N582, N605, N606, N607, N608, N609,
         N610, N611, N6120, N613, N614, N615, N616, N617, N618, N619, N620,
         N623, N624, N625, N626, N627, N628, N629, N630, N631, N632, N633,
         N634, N635, N636, N637, N638, N639, N640, N641, N642, N643, N644,
         N645, N646, N647, N648, N649, N650, N651, N652, N653, N654, N655,
         N656, N657, N658, N659, N660, N661, N662, N663, N664, N665, N666,
         N667, N668, N669, N670, N671, N672, N673, N674, N675, N676, N677,
         N678, N679, N680, N681, N682, N683, N684, N685, N686, N687, N688,
         N689, N690, N691, N692, N693, N694, N695, N696, N697, N698, N699,
         N700, N701, N702, N817, N821, N822, N823, N824, N825, N873, N874,
         N936, N937, N938, N939, N940, N941, N942, N943, N944, N945, N946,
         N947, N948, N949, N950, N951, N952, N953, N954, N955, N956, N957,
         N958, N959, N960, N961, N962, N963, N964, N965, N966, N967, N968,
         N969, N970, N971, N972, N973, N974, N975, N976, N977, N978, N979,
         N980, N981, N982, N983, N984, N985, N986, N987, N988, N989, N990,
         N991, N992, N993, N994, N995, N996, N997, N998, N999, N1000, N1001,
         N1002, N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011,
         N1012, N1013, N1014, N1015, N1016, SUB_X_283_4_N16, SUB_X_283_4_N15,
         SUB_X_283_4_N14, SUB_X_283_4_N13, SUB_X_283_4_N12, SUB_X_283_4_N11,
         SUB_X_283_4_N10, SUB_X_283_4_N9, SUB_X_283_4_N8, SUB_X_283_4_N7,
         SUB_X_283_4_N6, SUB_X_283_4_N5, SUB_X_283_4_N4, SUB_X_283_4_N3,
         SUB_X_283_4_N2, SUB_X_283_4_N1, ADD_X_283_3_N16, ADD_X_283_3_N15,
         ADD_X_283_3_N14, ADD_X_283_3_N13, ADD_X_283_3_N12, ADD_X_283_3_N11,
         ADD_X_283_3_N10, ADD_X_283_3_N9, ADD_X_283_3_N8, ADD_X_283_3_N7,
         ADD_X_283_3_N6, ADD_X_283_3_N5, ADD_X_283_3_N4, ADD_X_283_3_N3,
         ADD_X_283_3_N2, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12,
         N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26,
         N27, N119, N120, N121, N123, N124, N125, N126, N127, N128, N129, N130,
         N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, N141,
         N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152,
         N153, N155, N156, N157, N158, N159, N160, N161, N1620, N1630, N1640,
         N165, N166, N167, N168, N169, N170, N171, N172, N173, N174, N175,
         N176, N177, N178, N179, N180, N181, N182, N183, N184, N185, N186,
         N187, N188, N189, N190, N191, N192, N193, N194, N202, N203, N204,
         N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215,
         N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226,
         N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237,
         N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248,
         N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259,
         N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270,
         N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281,
         N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292,
         N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303,
         N304, N305, N306, N307, N308, N309, N310, N311, N312, N313, N314,
         N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325,
         N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336,
         N337, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347,
         N348, N349, N350, N351, N352, N353, N354, N355, N356, N357, N358,
         N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, N369,
         N370, N371, N372, N373, N374, N375, N376, N377, N378, N379, N380,
         N381, N382, N383, N384, N385, N386, N387, N388, N389, N390, N391,
         N392, N393, N394, N395, N396, N397, N398, N399, N400, N401, N402,
         N403, N404, N405, N406, N407, N408, N409, N410, N411, N413, N419,
         N422, N425, N426, N427, N428, N430, N433, N434, N435, N436, N437,
         N438, N439, N440, N441, N459, N489, N490, N491, N5000, N5010, N5020,
         N5050, N5080, N5110, N5140, N517, N520, N523, N526, N529, N532, N535,
         N538, N541, N544, N546, N547, N548, N549, N550, N551, N552, N553,
         N554, N555, N556, N557, N559, N560, N561, N563, N565, N566, N567,
         N568, N569, N570, N571, N572, N573, N574, N575, N576, N577, N578,
         N580, N581, N583, N5840, N5850, N586, N587, N588, N589, N590, N591,
         N592, N593, N594, N595, N596, N597, N598, N599, N600, N601, N602,
         N603, N604, N621, N622, N703, N704, N705, N706, N707, N708, N709,
         N710, N711, N712, N713, N714, N715, N716, N717, N718, N719, N720,
         N721, N722, N723, N724, N725, N726, N727, N728, N729, N730, N731,
         N732, N733, N734, N735, N736, N737, N738, N739, N740, N741, N742,
         N743, N744, N745, N746, N747, N748, N749, N750, N751, N752, N753,
         N754, N755, N756, N757, N758, N759, N760, N761, N762, N763, N764,
         N765, N766, N767, N768, N769, N770, N771, N772, N773, N774, N775,
         N776, N777, N778, N779, N780, N781, N782, N783, N784, N785, N786,
         N787, N788, N789, N790, N791, N792, N793, N794, N795, N796, N797,
         N798, N799, N800, N801, N802, N803, N804, N805, N806, N807, N808,
         N809, N810, N811, N812, N813, N814, N815, N816, N818, N819, N820,
         N826, N827, N828, N829, N830, N831, N832, N833, N834, N835, N836,
         N837, N838, N839, N840, N841, N842, N843, N844, N845, N846, N847,
         N848, N849, N850, N851, N852, N853, N854, N855, N856, N857, N858,
         N859, N860, N861, N862, N863, N864, N865, N866, N867, N868, N869,
         N870, N871, N872, N875, N876, N877, N878, N879, N880, N881, N882,
         N883, N884, N885, N886, N887, N888, N889, N890, N891, N892, N893,
         N894, N895, N896, N897, N898, N899, N900, N901, N902, N903, N904,
         N905, N906, N907, N908, N909, N910, N911, N912, N913, N914, N915,
         N916, N917, N918, N919, N920, N921, N922, N923, N924, N925, N926,
         N927, N928, N929, N930, N931, N932, N933, N934, N935, N1017, N1018,
         N1019, N1020, N1021, N1022, N1023, N1024, N1025, N1026, N1027, N1028,
         N1029, N1030, N1031, N1032, N1033, N1034, N1035, N1036, N1037, N1038,
         N1039, N1040, N1041, N1042, N1043, N1044, N1045, N1046, N1047, N1048,
         N1049, N1050, N1051, N1052, N1053, N1054, N1055, N1056, N1057, N1058,
         N1059, N1060, N1061, N1062, N1063, N1064, N1065, N1066, N1067, N1068,
         N1069, N1070, N1071, N1072, N1073, N1074, N1075, N1076, N1077, N1078,
         N1079, N1080, N1081, N1082, N1083, N1084, N1085, N1086, N1087, N1088,
         N1089, N1090, N1091, N1092, N1093, N1094, N1095, N1096, N1097, N1098,
         N1099, N1100, N1101, N1102, N1103, N1104, N1105, N1106, N1107, N1108,
         N1109, N1110, N1111, N1112, N1113, N1114, N1115, N1116, N1117, N1118,
         N1119, N1120, N1121, N1122, N1123, N1124, N1125, N1126, N1127, N1128,
         N1129, N1130, N1131, N1132, N1133, N1134, N1135, N1136, N1137, N1138,
         N1139, N11400, N1141, N1142, N1143, N1144, N1145, N1146, N1147, N1148,
         N1149, N1150, N1151, N1152, N1153, N1154, N1155, N1156, N1157, N1158,
         N1159, N1160, N1161, N1162, N1163, N1164, N1165, N1166, N1167, N1168,
         N1169, N1170, N1171, N1172, N1173, N1174, N1175;
  wire   [4:2] CODE_TYPE;
  wire   [2:0] OPER3_R3;
  wire   [1:0] STATE;
  wire   [2:0] NEXT_STATE;
  wire   [15:0] REG_A;
  wire   [15:0] REG_B;

  DFFSX2TF \pc_reg[2]  ( .D(N824), .CK(CLK), .SN(RST_N), .Q(N243), .QN(
        I_ADDR[3]) );
  DFFSX2TF \pc_reg[7]  ( .D(N873), .CK(CLK), .SN(RST_N), .Q(N233), .QN(
        I_ADDR[8]) );
  DFFSX2TF \pc_reg[5]  ( .D(N821), .CK(CLK), .SN(RST_N), .Q(N232), .QN(
        I_ADDR[6]) );
  DFFSX2TF \pc_reg[3]  ( .D(N823), .CK(CLK), .SN(RST_N), .Q(N231), .QN(
        I_ADDR[4]) );
  DFFSX2TF \state_reg[3]  ( .D(N558), .CK(CLK), .SN(RST_N), .Q(N562), .QN(N226) );
  TLATXLTF cf_buf_reg ( .G(N584), .D(N585), .Q(CF_BUF) );
  TLATXLTF \nxt_reg[0]  ( .G(N162), .D(N163), .Q(NXT[0]) );
  TLATXLTF \nxt_reg[1]  ( .G(N162), .D(N164), .Q(NXT[1]) );
  DFFSX2TF \pc_reg[6]  ( .D(N817), .CK(CLK), .SN(RST_N), .QN(I_ADDR[7]) );
  DFFSX2TF \pc_reg[4]  ( .D(N822), .CK(CLK), .SN(RST_N), .QN(I_ADDR[5]) );
  DFFSX2TF \pc_reg[1]  ( .D(N825), .CK(CLK), .SN(RST_N), .QN(I_ADDR[2]) );
  DFFSX2TF \pc_reg[0]  ( .D(N874), .CK(CLK), .SN(RST_N), .QN(I_ADDR[1]) );
  CMPR32X2TF \sub_x_283_4/U14  ( .A(N182), .B(REG_A[3]), .C(SUB_X_283_4_N14), 
        .CO(SUB_X_283_4_N13), .S(N503) );
  CMPR32X2TF \sub_x_283_4/U13  ( .A(N183), .B(REG_A[4]), .C(SUB_X_283_4_N13), 
        .CO(SUB_X_283_4_N12), .S(N504) );
  CMPR32X2TF \sub_x_283_4/U10  ( .A(N186), .B(REG_A[7]), .C(SUB_X_283_4_N10), 
        .CO(SUB_X_283_4_N9), .S(N507) );
  CMPR32X2TF \sub_x_283_4/U12  ( .A(N184), .B(REG_A[5]), .C(SUB_X_283_4_N12), 
        .CO(SUB_X_283_4_N11), .S(N505) );
  CMPR32X2TF \sub_x_283_4/U16  ( .A(N180), .B(REG_A[1]), .C(SUB_X_283_4_N16), 
        .CO(SUB_X_283_4_N15), .S(N501) );
  CMPR32X2TF \sub_x_283_4/U15  ( .A(N181), .B(REG_A[2]), .C(SUB_X_283_4_N15), 
        .CO(SUB_X_283_4_N14), .S(N502) );
  CMPR32X2TF \add_x_283_3/U12  ( .A(REG_A[5]), .B(REG_B[5]), .C(
        ADD_X_283_3_N12), .CO(ADD_X_283_3_N11), .S(N471) );
  CMPR32X2TF \add_x_283_3/U11  ( .A(REG_A[6]), .B(REG_B[6]), .C(
        ADD_X_283_3_N11), .CO(ADD_X_283_3_N10), .S(N472) );
  CMPR32X2TF \add_x_283_3/U10  ( .A(REG_A[7]), .B(REG_B[7]), .C(
        ADD_X_283_3_N10), .CO(ADD_X_283_3_N9), .S(N473) );
  CMPR32X2TF \add_x_283_3/U3  ( .A(REG_A[14]), .B(REG_B[14]), .C(
        ADD_X_283_3_N3), .CO(ADD_X_283_3_N2), .S(N480) );
  DFFNSRX2TF lowest_bit_reg ( .D(N1016), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        N123), .QN(N121) );
  DFFNSRXLTF \reg_C_reg[9]  ( .D(N518), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N424) );
  DFFNSRXLTF \reg_C_reg[11]  ( .D(N533), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N418) );
  DFFNSRXLTF \reg_C_reg[8]  ( .D(N5090), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N429) );
  DFFNSRXLTF \reg_C_reg[12]  ( .D(N524), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N423) );
  DFFNSRXLTF \reg_C_reg[10]  ( .D(N527), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N421) );
  DFFNSRXLTF \reg_C_reg[13]  ( .D(N530), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N420) );
  DFFNSRXLTF \reg_C_reg[14]  ( .D(N536), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N417) );
  DFFNSRXLTF \reg_C_reg[15]  ( .D(N542), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N412) );
  DFFNSRXLTF is_i_addr_reg ( .D(N114), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        IS_I_ADDR) );
  DFFNSRXLTF dw_reg ( .D(N612), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(D_WE) );
  DFFRX4TF \reg_A_reg[0]  ( .D(N464), .CK(CLK), .RN(RST_N), .Q(REG_A[0]), .QN(
        N206) );
  DFFRX4TF \reg_B_reg[2]  ( .D(N519), .CK(CLK), .RN(RST_N), .Q(REG_B[2]), .QN(
        N181) );
  DFFRX4TF \reg_B_reg[1]  ( .D(N537), .CK(CLK), .RN(RST_N), .Q(REG_B[1]), .QN(
        N180) );
  DFFRX4TF \reg_B_reg[0]  ( .D(N543), .CK(CLK), .RN(RST_N), .Q(REG_B[0]), .QN(
        N1150) );
  DFFRX1TF \smdr_reg[0]  ( .D(N488), .CK(CLK), .RN(RST_N), .QN(N620) );
  DFFRX1TF \smdr_reg[13]  ( .D(N4760), .CK(CLK), .RN(RST_N), .QN(N607) );
  DFFRX1TF \smdr_reg[10]  ( .D(N4790), .CK(CLK), .RN(RST_N), .QN(N610) );
  DFFRX1TF \smdr_reg[8]  ( .D(N4810), .CK(CLK), .RN(RST_N), .QN(N6120) );
  DFFRX1TF \smdr_reg[14]  ( .D(N4750), .CK(CLK), .RN(RST_N), .QN(N606) );
  DFFRX1TF \smdr_reg[12]  ( .D(N4770), .CK(CLK), .RN(RST_N), .QN(N608) );
  DFFRX1TF \smdr_reg[7]  ( .D(N462), .CK(CLK), .RN(RST_N), .QN(N613) );
  DFFRX1TF \smdr_reg[3]  ( .D(N458), .CK(CLK), .RN(RST_N), .QN(N617) );
  DFFRX1TF \smdr_reg[11]  ( .D(N4780), .CK(CLK), .RN(RST_N), .QN(N609) );
  DFFRX1TF \smdr_reg[2]  ( .D(N486), .CK(CLK), .RN(RST_N), .QN(N618) );
  DFFRX1TF \smdr_reg[6]  ( .D(N483), .CK(CLK), .RN(RST_N), .QN(N614) );
  DFFRX1TF \smdr_reg[4]  ( .D(N485), .CK(CLK), .RN(RST_N), .QN(N616) );
  DFFRX1TF \smdr_reg[15]  ( .D(N4820), .CK(CLK), .RN(RST_N), .QN(N605) );
  DFFRX1TF \smdr_reg[9]  ( .D(N4800), .CK(CLK), .RN(RST_N), .QN(N611) );
  DFFRX1TF \smdr_reg[5]  ( .D(N484), .CK(CLK), .RN(RST_N), .QN(N615) );
  DFFRX1TF \smdr_reg[1]  ( .D(N487), .CK(CLK), .RN(RST_N), .QN(N619) );
  DFFRX1TF \id_ir_reg[7]  ( .D(N463), .CK(CLK), .RN(RST_N), .QN(N432) );
  DFFRX1TF \id_ir_reg[3]  ( .D(N4700), .CK(CLK), .RN(RST_N), .QN(N431) );
  DFFRX1TF \id_ir_reg[9]  ( .D(N498), .CK(CLK), .RN(RST_N), .Q(N124), .QN(N25)
         );
  DFFRX1TF \gr_reg[2][14]  ( .D(N952), .CK(CLK), .RN(RST_N), .QN(N656) );
  DFFRX1TF \gr_reg[2][13]  ( .D(N953), .CK(CLK), .RN(RST_N), .QN(N657) );
  DFFRX1TF \gr_reg[2][15]  ( .D(N951), .CK(CLK), .RN(RST_N), .QN(N655) );
  DFFRX1TF \gr_reg[4][14]  ( .D(N936), .CK(CLK), .RN(RST_N), .QN(N624) );
  DFFRX1TF \gr_reg[4][13]  ( .D(N937), .CK(CLK), .RN(RST_N), .QN(N625) );
  DFFRX1TF \gr_reg[4][12]  ( .D(N938), .CK(CLK), .RN(RST_N), .QN(N626) );
  DFFRX1TF \gr_reg[4][11]  ( .D(N939), .CK(CLK), .RN(RST_N), .QN(N627) );
  DFFRX1TF \gr_reg[4][10]  ( .D(N940), .CK(CLK), .RN(RST_N), .QN(N628) );
  DFFRX1TF \gr_reg[4][15]  ( .D(N1015), .CK(CLK), .RN(RST_N), .QN(N623) );
  DFFRX1TF \gr_reg[1][15]  ( .D(N959), .CK(CLK), .RN(RST_N), .QN(N671) );
  DFFRX1TF \gr_reg[1][14]  ( .D(N960), .CK(CLK), .RN(RST_N), .QN(N672) );
  DFFRX1TF \gr_reg[1][13]  ( .D(N961), .CK(CLK), .RN(RST_N), .QN(N673) );
  DFFRX1TF \gr_reg[1][12]  ( .D(N962), .CK(CLK), .RN(RST_N), .QN(N674) );
  DFFRX1TF \gr_reg[1][11]  ( .D(N963), .CK(CLK), .RN(RST_N), .QN(N675) );
  DFFRX1TF \gr_reg[1][10]  ( .D(N964), .CK(CLK), .RN(RST_N), .QN(N676) );
  DFFRX1TF \gr_reg[1][9]  ( .D(N965), .CK(CLK), .RN(RST_N), .QN(N677) );
  DFFRX1TF \gr_reg[1][8]  ( .D(N966), .CK(CLK), .RN(RST_N), .QN(N678) );
  DFFRX1TF \gr_reg[0][15]  ( .D(N967), .CK(CLK), .RN(RST_N), .QN(N687) );
  DFFRX1TF \gr_reg[0][14]  ( .D(N968), .CK(CLK), .RN(RST_N), .QN(N688) );
  DFFRX1TF \gr_reg[0][13]  ( .D(N969), .CK(CLK), .RN(RST_N), .QN(N689) );
  DFFRX1TF \gr_reg[0][12]  ( .D(N970), .CK(CLK), .RN(RST_N), .QN(N690) );
  DFFRX1TF \gr_reg[0][11]  ( .D(N971), .CK(CLK), .RN(RST_N), .QN(N691) );
  DFFRX1TF \gr_reg[0][10]  ( .D(N972), .CK(CLK), .RN(RST_N), .QN(N692) );
  DFFRX1TF \gr_reg[0][9]  ( .D(N973), .CK(CLK), .RN(RST_N), .QN(N693) );
  DFFRX1TF \gr_reg[0][8]  ( .D(N974), .CK(CLK), .RN(RST_N), .QN(N694) );
  DFFRX1TF \gr_reg[1][7]  ( .D(N999), .CK(CLK), .RN(RST_N), .QN(N679) );
  DFFRX1TF \gr_reg[1][6]  ( .D(N1000), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[6]), 
        .QN(N680) );
  DFFRX1TF \gr_reg[0][5]  ( .D(N1009), .CK(CLK), .RN(RST_N), .QN(N697) );
  DFFRX1TF \gr_reg[0][3]  ( .D(N1011), .CK(CLK), .RN(RST_N), .QN(N699) );
  DFFRX1TF \gr_reg[0][7]  ( .D(N1007), .CK(CLK), .RN(RST_N), .QN(N695) );
  DFFRX1TF \gr_reg[0][6]  ( .D(N1008), .CK(CLK), .RN(RST_N), .QN(N696) );
  DFFRX1TF \gr_reg[0][4]  ( .D(N1010), .CK(CLK), .RN(RST_N), .QN(N698) );
  DFFRX1TF \gr_reg[0][2]  ( .D(N1012), .CK(CLK), .RN(RST_N), .QN(N700) );
  DFFRX1TF \gr_reg[0][1]  ( .D(N1013), .CK(CLK), .RN(RST_N), .QN(N701) );
  DFFRX1TF \gr_reg[0][0]  ( .D(N1014), .CK(CLK), .RN(RST_N), .QN(N702) );
  DFFRX2TF \state_reg[2]  ( .D(NEXT_STATE[2]), .CK(CLK), .RN(RST_N), .Q(N230), 
        .QN(N564) );
  DFFRX2TF \reg_A_reg[14]  ( .D(N534), .CK(CLK), .RN(RST_N), .Q(REG_A[14]), 
        .QN(N204) );
  DFFRX2TF \reg_A_reg[13]  ( .D(N528), .CK(CLK), .RN(RST_N), .Q(REG_A[13]), 
        .QN(N211) );
  DFFRX2TF \reg_A_reg[11]  ( .D(N531), .CK(CLK), .RN(RST_N), .Q(REG_A[11]), 
        .QN(N220) );
  DFFRX2TF \reg_A_reg[10]  ( .D(N525), .CK(CLK), .RN(RST_N), .Q(REG_A[10]), 
        .QN(N214) );
  DFFRX2TF \reg_A_reg[9]  ( .D(N5160), .CK(CLK), .RN(RST_N), .Q(REG_A[9]), 
        .QN(N213) );
  DFFRX2TF \reg_A_reg[8]  ( .D(N5070), .CK(CLK), .RN(RST_N), .Q(REG_A[8]), 
        .QN(N215) );
  DFFRX2TF \reg_A_reg[5]  ( .D(N5040), .CK(CLK), .RN(RST_N), .Q(REG_A[5]), 
        .QN(N217) );
  DFFRX2TF \reg_A_reg[1]  ( .D(N465), .CK(CLK), .RN(RST_N), .Q(REG_A[1]), .QN(
        N202) );
  DFFRX2TF \state_reg[0]  ( .D(NEXT_STATE[0]), .CK(CLK), .RN(RST_N), .Q(
        STATE[0]), .QN(N207) );
  DFFRX2TF \reg_A_reg[15]  ( .D(N540), .CK(CLK), .RN(RST_N), .Q(REG_A[15]), 
        .QN(N210) );
  DFFRX2TF \reg_A_reg[7]  ( .D(N461), .CK(CLK), .RN(RST_N), .Q(REG_A[7]), .QN(
        N218) );
  DFFRX2TF \reg_A_reg[2]  ( .D(N4660), .CK(CLK), .RN(RST_N), .Q(REG_A[2]), 
        .QN(N219) );
  DFFRX2TF \reg_A_reg[12]  ( .D(N522), .CK(CLK), .RN(RST_N), .Q(REG_A[12]), 
        .QN(N216) );
  DFFRX2TF \reg_A_reg[3]  ( .D(N457), .CK(CLK), .RN(RST_N), .Q(REG_A[3]), .QN(
        N221) );
  DFFRX2TF \reg_A_reg[4]  ( .D(N5130), .CK(CLK), .RN(RST_N), .Q(REG_A[4]), 
        .QN(N209) );
  DFFRX2TF \reg_A_reg[6]  ( .D(N5100), .CK(CLK), .RN(RST_N), .Q(REG_A[6]), 
        .QN(N212) );
  DFFRX2TF \reg_B_reg[13]  ( .D(N446), .CK(CLK), .RN(RST_N), .Q(REG_B[13]), 
        .QN(N192) );
  DFFRX2TF \reg_B_reg[12]  ( .D(N449), .CK(CLK), .RN(RST_N), .Q(REG_B[12]), 
        .QN(N191) );
  DFFRX2TF \reg_B_reg[15]  ( .D(N443), .CK(CLK), .RN(RST_N), .Q(REG_B[15]), 
        .QN(N194) );
  DFFRX2TF \reg_B_reg[11]  ( .D(N445), .CK(CLK), .RN(RST_N), .Q(REG_B[11]), 
        .QN(N190) );
  DFFRX2TF \reg_B_reg[9]  ( .D(N450), .CK(CLK), .RN(RST_N), .Q(REG_B[9]), .QN(
        N188) );
  DFFRX2TF nf_reg ( .D(N442), .CK(CLK), .RN(RST_N), .Q(NF), .QN(N234) );
  DFFRX2TF \reg_B_reg[7]  ( .D(N455), .CK(CLK), .RN(RST_N), .Q(REG_B[7]), .QN(
        N186) );
  DFFRX2TF \reg_B_reg[3]  ( .D(N456), .CK(CLK), .RN(RST_N), .Q(REG_B[3]), .QN(
        N182) );
  DFFRX2TF \reg_B_reg[6]  ( .D(N452), .CK(CLK), .RN(RST_N), .Q(REG_B[6]), .QN(
        N185) );
  DFFRX2TF \reg_B_reg[5]  ( .D(N454), .CK(CLK), .RN(RST_N), .Q(REG_B[5]), .QN(
        N184) );
  DFFRX2TF \reg_B_reg[4]  ( .D(N451), .CK(CLK), .RN(RST_N), .Q(REG_B[4]), .QN(
        N183) );
  DFFRX2TF \reg_B_reg[10]  ( .D(N447), .CK(CLK), .RN(RST_N), .Q(REG_B[10]), 
        .QN(N189) );
  DFFRX2TF \reg_B_reg[8]  ( .D(N453), .CK(CLK), .RN(RST_N), .Q(REG_B[8]), .QN(
        N187) );
  DFFRX2TF \reg_B_reg[14]  ( .D(N444), .CK(CLK), .RN(RST_N), .Q(REG_B[14]), 
        .QN(N193) );
  DFFRX2TF zf_reg ( .D(N448), .CK(CLK), .RN(RST_N), .Q(ZF), .QN(N235) );
  DFFRX2TF \id_ir_reg[6]  ( .D(N4670), .CK(CLK), .RN(RST_N), .Q(N236), .QN(
        N414) );
  DFFRX2TF \id_ir_reg[5]  ( .D(N4680), .CK(CLK), .RN(RST_N), .Q(N237), .QN(
        N415) );
  DFFRX2TF \id_ir_reg[4]  ( .D(N4690), .CK(CLK), .RN(RST_N), .Q(N238), .QN(
        N416) );
  DFFRX2TF \id_ir_reg[2]  ( .D(N4710), .CK(CLK), .RN(RST_N), .Q(OPER3_R3[2]), 
        .QN(N239) );
  DFFRX2TF \id_ir_reg[0]  ( .D(N4730), .CK(CLK), .RN(RST_N), .Q(OPER3_R3[0]), 
        .QN(N228) );
  DFFRX2TF \id_ir_reg[14]  ( .D(N493), .CK(CLK), .RN(RST_N), .Q(CODE_TYPE[3]), 
        .QN(N229) );
  DFFRX2TF \id_ir_reg[13]  ( .D(N494), .CK(CLK), .RN(RST_N), .Q(CODE_TYPE[2]), 
        .QN(N225) );
  DFFRX2TF \id_ir_reg[12]  ( .D(N495), .CK(CLK), .RN(RST_N), .Q(N208), .QN(N26) );
  DFFRX2TF \id_ir_reg[10]  ( .D(N497), .CK(CLK), .RN(RST_N), .Q(\OPER1_R1[2] ), 
        .QN(N227) );
  DFFRX2TF \id_ir_reg[8]  ( .D(N499), .CK(CLK), .RN(RST_N), .Q(N222), .QN(N582) );
  DFFRX2TF \id_ir_reg[15]  ( .D(N492), .CK(CLK), .RN(RST_N), .Q(CODE_TYPE[4]), 
        .QN(N205) );
  DFFRX2TF \id_ir_reg[11]  ( .D(N496), .CK(CLK), .RN(RST_N), .Q(N203), .QN(
        N579) );
  DFFRX2TF \id_ir_reg[1]  ( .D(N4720), .CK(CLK), .RN(RST_N), .Q(OPER3_R3[1]), 
        .QN(N223) );
  DFFRX2TF \gr_reg[3][14]  ( .D(N944), .CK(CLK), .RN(RST_N), .Q(N241), .QN(
        N640) );
  DFFRX2TF \gr_reg[3][13]  ( .D(N945), .CK(CLK), .RN(RST_N), .Q(N240), .QN(
        N641) );
  DFFRX2TF \gr_reg[3][12]  ( .D(N946), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTB[12]), .QN(N642) );
  DFFRX2TF \gr_reg[3][11]  ( .D(N947), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTB[11]), .QN(N643) );
  DFFRX2TF \gr_reg[3][10]  ( .D(N948), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTB[10]), .QN(N644) );
  DFFRX2TF \gr_reg[3][9]  ( .D(N949), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[9]), 
        .QN(N645) );
  DFFRX2TF \gr_reg[3][8]  ( .D(N950), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[8]), 
        .QN(N646) );
  DFFRX2TF \gr_reg[2][12]  ( .D(N954), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTA[12]), .QN(N658) );
  DFFRX2TF \gr_reg[2][11]  ( .D(N955), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTA[11]), .QN(N659) );
  DFFRX2TF \gr_reg[2][10]  ( .D(N956), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTA[10]), .QN(N660) );
  DFFRX2TF \gr_reg[2][9]  ( .D(N957), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[9]), 
        .QN(N661) );
  DFFRX2TF \gr_reg[2][8]  ( .D(N958), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[8]), 
        .QN(N662) );
  DFFRX2TF \gr_reg[3][15]  ( .D(N943), .CK(CLK), .RN(RST_N), .Q(N242), .QN(
        N639) );
  DFFRX2TF \gr_reg[4][9]  ( .D(N941), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[9]), 
        .QN(N629) );
  DFFRX2TF \gr_reg[4][8]  ( .D(N942), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[8]), 
        .QN(N630) );
  DFFRX2TF \gr_reg[4][5]  ( .D(N977), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[5]), 
        .QN(N633) );
  DFFRX2TF \gr_reg[4][3]  ( .D(N979), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[3]), 
        .QN(N635) );
  DFFRX2TF \gr_reg[4][7]  ( .D(N975), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[7]), 
        .QN(N631) );
  DFFRX2TF \gr_reg[4][6]  ( .D(N976), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[6]), 
        .QN(N632) );
  DFFRX2TF \gr_reg[4][4]  ( .D(N978), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[4]), 
        .QN(N634) );
  DFFRX2TF \gr_reg[4][2]  ( .D(N980), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[2]), 
        .QN(N636) );
  DFFRX2TF \gr_reg[4][1]  ( .D(N981), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[1]), 
        .QN(N637) );
  DFFRX2TF \gr_reg[4][0]  ( .D(N982), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[0]), 
        .QN(N638) );
  DFFRX2TF \gr_reg[3][5]  ( .D(N985), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[5]), 
        .QN(N649) );
  DFFRX2TF \gr_reg[3][3]  ( .D(N987), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[3]), 
        .QN(N651) );
  DFFRX2TF \gr_reg[2][5]  ( .D(N993), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[5]), 
        .QN(N665) );
  DFFRX2TF \gr_reg[2][3]  ( .D(N995), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[3]), 
        .QN(N667) );
  DFFRX2TF \gr_reg[3][7]  ( .D(N983), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[7]), 
        .QN(N647) );
  DFFRX2TF \gr_reg[3][6]  ( .D(N984), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[6]), 
        .QN(N648) );
  DFFRX2TF \gr_reg[3][4]  ( .D(N986), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[4]), 
        .QN(N650) );
  DFFRX2TF \gr_reg[3][2]  ( .D(N988), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[2]), 
        .QN(N652) );
  DFFRX2TF \gr_reg[3][1]  ( .D(N989), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[1]), 
        .QN(N653) );
  DFFRX2TF \gr_reg[3][0]  ( .D(N990), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[0]), 
        .QN(N654) );
  DFFRX2TF \gr_reg[2][7]  ( .D(N991), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[7]), 
        .QN(N663) );
  DFFRX2TF \gr_reg[2][6]  ( .D(N992), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[6]), 
        .QN(N664) );
  DFFRX2TF \gr_reg[2][4]  ( .D(N994), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[4]), 
        .QN(N666) );
  DFFRX2TF \gr_reg[2][2]  ( .D(N996), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[2]), 
        .QN(N668) );
  DFFRX2TF \gr_reg[2][1]  ( .D(N997), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[1]), 
        .QN(N669) );
  DFFRX2TF \gr_reg[2][0]  ( .D(N998), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[0]), 
        .QN(N670) );
  DFFRX2TF \gr_reg[1][5]  ( .D(N1001), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[5]), 
        .QN(N681) );
  DFFRX2TF \gr_reg[1][3]  ( .D(N1003), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[3]), 
        .QN(N683) );
  DFFRX2TF \gr_reg[1][4]  ( .D(N1002), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[4]), 
        .QN(N682) );
  DFFRX2TF \gr_reg[1][2]  ( .D(N1004), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[2]), 
        .QN(N684) );
  DFFRX2TF \gr_reg[1][1]  ( .D(N1005), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[1]), 
        .QN(N685) );
  DFFRX2TF \gr_reg[1][0]  ( .D(N1006), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[0]), 
        .QN(N686) );
  DFFRX1TF \state_reg[1]  ( .D(NEXT_STATE[1]), .CK(CLK), .RN(RST_N), .Q(
        STATE[1]) );
  DFFRX1TF cf_reg ( .D(N4740), .CK(CLK), .RN(RST_N), .Q(CF) );
  DFFNSRX2TF \reg_C_reg[5]  ( .D(N5060), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[6]) );
  DFFNSRX2TF \reg_C_reg[3]  ( .D(N460), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[4]) );
  DFFNSRX2TF \reg_C_reg[0]  ( .D(N545), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[1]) );
  DFFNSRX2TF \reg_C_reg[7]  ( .D(N5030), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[8]) );
  DFFNSRX2TF \reg_C_reg[2]  ( .D(N521), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[3]) );
  DFFNSRX2TF \reg_C_reg[6]  ( .D(N5120), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[7]) );
  DFFNSRX2TF \reg_C_reg[4]  ( .D(N5150), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[5]) );
  DFFNSRX2TF \reg_C_reg[1]  ( .D(N539), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[2]) );
  OR3X1TF U3 ( .A(N26), .B(N860), .C(N358), .Y(N791) );
  INVX2TF U4 ( .A(N590), .Y(N748) );
  ADDFX2TF U5 ( .A(N192), .B(REG_A[13]), .CI(SUB_X_283_4_N4), .CO(
        SUB_X_283_4_N3), .S(N513) );
  AOI21X1TF U6 ( .A0(N479), .A1(N148), .B0(N759), .Y(N761) );
  NAND3X1TF U7 ( .A(N26), .B(N893), .C(N859), .Y(N782) );
  NAND2X1TF U8 ( .A(N562), .B(N207), .Y(N345) );
  NAND2X1TF U9 ( .A(N130), .B(N890), .Y(N1141) );
  AOI211X2TF U10 ( .A0(N798), .A1(N719), .B0(N402), .C0(N401), .Y(N1166) );
  CLKBUFX2TF U11 ( .A(N1159), .Y(N169) );
  ADDFX2TF U12 ( .A(REG_A[15]), .B(REG_B[15]), .CI(ADD_X_283_3_N2), .CO(N482), 
        .S(N481) );
  AOI211X1TF U13 ( .A0(REG_A[10]), .A1(N173), .B0(N604), .C0(N567), .Y(N1) );
  NAND2X1TF U14 ( .A(N5000), .B(N1), .Y(N406) );
  AOI21X1TF U15 ( .A0(N153), .A1(REG_A[4]), .B0(N603), .Y(N2) );
  NAND3X1TF U16 ( .A(N491), .B(N740), .C(N2), .Y(N719) );
  OA21XLTF U17 ( .A0(I_ADDR[1]), .A1(I_ADDR[2]), .B0(N317), .Y(N3) );
  AOI222XLTF U18 ( .A0(I_ADDR[2]), .A1(N331), .B0(D_ADDR[2]), .B1(N330), .C0(
        N328), .C1(N3), .Y(N825) );
  NOR4XLTF U19 ( .A(N1169), .B(N1160), .C(N1164), .D(N1067), .Y(N4) );
  NOR4XLTF U20 ( .A(N1081), .B(N1061), .C(N1055), .D(N1074), .Y(N5) );
  NOR3X1TF U21 ( .A(N1089), .B(N1118), .C(N1088), .Y(N6) );
  NAND4X1TF U22 ( .A(N4), .B(N5), .C(N6), .D(N1096), .Y(N7) );
  NAND4BX1TF U23 ( .AN(N918), .B(N1132), .C(N1166), .D(N1142), .Y(N8) );
  OAI2BB2XLTF U24 ( .B0(N7), .B1(N8), .A0N(N918), .A1N(ZF), .Y(N448) );
  OA22X1TF U25 ( .A0(N334), .A1(N333), .B0(N343), .B1(N336), .Y(N9) );
  NAND2X1TF U26 ( .A(N906), .B(START), .Y(N10) );
  OA22X1TF U27 ( .A0(N340), .A1(N337), .B0(STATE[1]), .B1(N10), .Y(N11) );
  NAND4X1TF U28 ( .A(N1144), .B(N344), .C(N9), .D(N11), .Y(NEXT_STATE[0]) );
  OA21XLTF U29 ( .A0(N321), .A1(I_ADDR[5]), .B0(N324), .Y(N12) );
  AOI222XLTF U30 ( .A0(I_ADDR[5]), .A1(N331), .B0(D_ADDR[5]), .B1(N330), .C0(
        N328), .C1(N12), .Y(N822) );
  CLKINVX1TF U31 ( .A(N893), .Y(N13) );
  OAI21X1TF U32 ( .A0(N208), .A1(N579), .B0(N13), .Y(N14) );
  AOI211X1TF U33 ( .A0(N349), .A1(CODE_TYPE[2]), .B0(N852), .C0(CODE_TYPE[3]), 
        .Y(N15) );
  OAI21X1TF U34 ( .A0(N26), .A1(N354), .B0(N350), .Y(N16) );
  AOI211X1TF U35 ( .A0(CODE_TYPE[4]), .A1(N14), .B0(N15), .C0(N16), .Y(N147)
         );
  OAI22X1TF U36 ( .A0(N1142), .A1(N1141), .B0(N1165), .B1(N1143), .Y(N17) );
  AOI21X1TF U37 ( .A0(IO_DATAINA[15]), .A1(N169), .B0(N17), .Y(N18) );
  OAI21X1TF U38 ( .A0(N131), .A1(N412), .B0(N18), .Y(N542) );
  OA21XLTF U39 ( .A0(N329), .A1(I_ADDR[7]), .B0(N327), .Y(N19) );
  AOI222XLTF U40 ( .A0(I_ADDR[7]), .A1(N331), .B0(D_ADDR[7]), .B1(N330), .C0(
        N328), .C1(N19), .Y(N817) );
  AOI21X1TF U41 ( .A0(N153), .A1(REG_A[11]), .B0(N422), .Y(N20) );
  NAND3X1TF U42 ( .A(N419), .B(N551), .C(N20), .Y(N731) );
  OAI22X1TF U43 ( .A0(N1142), .A1(N1143), .B0(N1162), .B1(N1141), .Y(N21) );
  AOI21X1TF U44 ( .A0(IO_DATAINA[14]), .A1(N169), .B0(N21), .Y(N22) );
  OAI21X1TF U45 ( .A0(N131), .A1(N417), .B0(N22), .Y(N536) );
  AOI21X1TF U46 ( .A0(N317), .A1(N243), .B0(N323), .Y(N23) );
  AOI222XLTF U47 ( .A0(I_ADDR[3]), .A1(N331), .B0(N23), .B1(N318), .C0(N330), 
        .C1(D_ADDR[3]), .Y(N824) );
  OR2X2TF U48 ( .A(REG_B[1]), .B(N1150), .Y(N24) );
  INVXLTF U49 ( .A(N26), .Y(N27) );
  NAND3X1TF U50 ( .A(N1175), .B(N1174), .C(N1173), .Y(N545) );
  NAND2XLTF U70 ( .A(N153), .B(REG_A[3]), .Y(N433) );
  NAND2XLTF U71 ( .A(N590), .B(N182), .Y(N396) );
  OR3X1TF U72 ( .A(REG_B[2]), .B(REG_B[3]), .C(N782), .Y(N805) );
  NAND2XLTF U73 ( .A(N173), .B(REG_A[11]), .Y(N352) );
  CMPR22X2TF U74 ( .A(REG_B[0]), .B(REG_A[0]), .CO(ADD_X_283_3_N16), .S(N466)
         );
  OR3X1TF U75 ( .A(N139), .B(N892), .C(N891), .Y(N1157) );
  AO22X1TF U76 ( .A0(\OPER1_R1[2] ), .A1(N870), .B0(N869), .B1(N236), .Y(N1137) );
  AO22X1TF U77 ( .A0(N886), .A1(N870), .B0(N416), .B1(N867), .Y(N1135) );
  NAND2XLTF U78 ( .A(N153), .B(REG_A[2]), .Y(N739) );
  OR4X2TF U79 ( .A(N26), .B(N882), .C(N881), .D(N880), .Y(N1042) );
  NAND3XLTF U80 ( .A(N336), .B(N344), .C(N335), .Y(NEXT_STATE[1]) );
  NAND3X2TF U81 ( .A(STATE[0]), .B(N365), .C(N226), .Y(N273) );
  INVX2TF U82 ( .A(N548), .Y(N119) );
  NAND2XLTF U83 ( .A(N548), .B(REG_A[6]), .Y(N549) );
  OR2X2TF U84 ( .A(REG_B[0]), .B(N1124), .Y(N752) );
  CLKINVX1TF U85 ( .A(N860), .Y(N348) );
  OR3X2TF U86 ( .A(N564), .B(STATE[1]), .C(N345), .Y(N1144) );
  NAND2BX2TF U87 ( .AN(REG_A[0]), .B(REG_B[0]), .Y(SUB_X_283_4_N16) );
  OAI31X2TF U88 ( .A0(REG_B[3]), .A1(N748), .A2(N716), .B0(N405), .Y(N410) );
  OAI21X1TF U89 ( .A0(N638), .A1(N172), .B0(N1155), .Y(N543) );
  OAI21XLTF U90 ( .A0(N680), .A1(N161), .B0(N1073), .Y(N5100) );
  OAI21X1TF U91 ( .A0(N627), .A1(N176), .B0(N932), .Y(N4780) );
  OAI21X1TF U92 ( .A0(N638), .A1(N175), .B0(N1048), .Y(N488) );
  OAI21X1TF U93 ( .A0(N628), .A1(N175), .B0(N935), .Y(N4790) );
  OAI21X1TF U94 ( .A0(N629), .A1(N176), .B0(N1019), .Y(N4800) );
  OAI21X1TF U95 ( .A0(N623), .A1(N176), .B0(N1025), .Y(N4820) );
  OAI21X1TF U96 ( .A0(N631), .A1(N172), .B0(N847), .Y(N455) );
  OAI21X1TF U97 ( .A0(N630), .A1(N175), .B0(N1022), .Y(N4810) );
  OAI21X1TF U98 ( .A0(N632), .A1(N176), .B0(N1028), .Y(N483) );
  OAI21X1TF U99 ( .A0(N634), .A1(N176), .B0(N1034), .Y(N485) );
  OAI21X1TF U100 ( .A0(N637), .A1(N172), .B0(N1128), .Y(N537) );
  OAI21X1TF U101 ( .A0(N625), .A1(N175), .B0(N926), .Y(N4760) );
  OAI21X1TF U102 ( .A0(N626), .A1(N176), .B0(N929), .Y(N4770) );
  OAI21X1TF U103 ( .A0(N637), .A1(N176), .B0(N1040), .Y(N487) );
  OAI21X1TF U104 ( .A0(N636), .A1(N172), .B0(N1095), .Y(N519) );
  OAI21X1TF U105 ( .A0(N624), .A1(N176), .B0(N923), .Y(N4750) );
  OAI21X1TF U106 ( .A0(N633), .A1(N176), .B0(N1031), .Y(N484) );
  OAI21X1TF U107 ( .A0(N636), .A1(N176), .B0(N1037), .Y(N486) );
  AOI211X1TF U108 ( .A0(N1047), .A1(IO_DATAOUTB[1]), .B0(N1039), .C0(N1038), 
        .Y(N1040) );
  AOI211X1TF U109 ( .A0(N1047), .A1(IO_DATAOUTB[12]), .B0(N928), .C0(N927), 
        .Y(N929) );
  AOI211X1TF U110 ( .A0(N1047), .A1(N240), .B0(N925), .C0(N924), .Y(N926) );
  AOI211X1TF U111 ( .A0(N167), .A1(IO_DATAOUTB[6]), .B0(N1027), .C0(N1026), 
        .Y(N1028) );
  AOI211X1TF U112 ( .A0(N167), .A1(IO_DATAOUTB[2]), .B0(N1036), .C0(N1035), 
        .Y(N1037) );
  AOI211X1TF U113 ( .A0(N1047), .A1(IO_DATAOUTB[5]), .B0(N1030), .C0(N1029), 
        .Y(N1031) );
  AOI211X1TF U114 ( .A0(N1047), .A1(N241), .B0(N922), .C0(N921), .Y(N923) );
  AOI211X1TF U115 ( .A0(N167), .A1(IO_DATAOUTB[4]), .B0(N1033), .C0(N1032), 
        .Y(N1034) );
  AOI211X1TF U116 ( .A0(N1047), .A1(IO_DATAOUTB[8]), .B0(N1021), .C0(N1020), 
        .Y(N1022) );
  AOI211X1TF U117 ( .A0(N1047), .A1(N242), .B0(N1024), .C0(N1023), .Y(N1025)
         );
  AOI211X1TF U118 ( .A0(N1047), .A1(IO_DATAOUTB[10]), .B0(N934), .C0(N933), 
        .Y(N935) );
  AOI211X1TF U119 ( .A0(N167), .A1(IO_DATAOUTB[11]), .B0(N931), .C0(N930), .Y(
        N932) );
  AOI211X1TF U120 ( .A0(N1047), .A1(IO_DATAOUTB[9]), .B0(N1018), .C0(N1017), 
        .Y(N1019) );
  OAI22X1TF U121 ( .A0(N690), .A1(N1044), .B0(N658), .B1(N150), .Y(N927) );
  OAI22X1TF U122 ( .A0(N688), .A1(N1044), .B0(N656), .B1(N150), .Y(N921) );
  AOI22X1TF U123 ( .A0(N278), .A1(N286), .B0(N685), .B1(N277), .Y(N1005) );
  AOI22X1TF U124 ( .A0(N303), .A1(N306), .B0(N655), .B1(N302), .Y(N951) );
  OAI22X1TF U125 ( .A0(N689), .A1(N1044), .B0(N657), .B1(N150), .Y(N924) );
  OAI22X1TF U126 ( .A0(N702), .A1(N1044), .B0(N670), .B1(N150), .Y(N1045) );
  OAI22X1TF U127 ( .A0(N694), .A1(N1044), .B0(N662), .B1(N150), .Y(N1020) );
  AOI22X1TF U128 ( .A0(N301), .A1(N315), .B0(N672), .B1(N300), .Y(N960) );
  OAI22X1TF U129 ( .A0(N692), .A1(N1044), .B0(N660), .B1(N150), .Y(N933) );
  AOI22X1TF U130 ( .A0(N301), .A1(N311), .B0(N675), .B1(N300), .Y(N963) );
  AOI22X1TF U131 ( .A0(N301), .A1(N308), .B0(N678), .B1(N300), .Y(N966) );
  AOI22X1TF U132 ( .A0(N307), .A1(N308), .B0(N646), .B1(N305), .Y(N950) );
  AOI22X1TF U133 ( .A0(N280), .A1(N290), .B0(N665), .B1(N279), .Y(N993) );
  AOI22X1TF U134 ( .A0(N283), .A1(N285), .B0(N654), .B1(N282), .Y(N990) );
  AOI22X1TF U135 ( .A0(N280), .A1(N288), .B0(N667), .B1(N279), .Y(N995) );
  AOI22X1TF U136 ( .A0(N307), .A1(N313), .B0(N641), .B1(N305), .Y(N945) );
  AOI22X1TF U137 ( .A0(N283), .A1(N286), .B0(N653), .B1(N282), .Y(N989) );
  AOI22X1TF U138 ( .A0(N283), .A1(N287), .B0(N652), .B1(N282), .Y(N988) );
  AOI22X1TF U139 ( .A0(N303), .A1(N309), .B0(N661), .B1(N302), .Y(N957) );
  AOI22X1TF U140 ( .A0(N307), .A1(N315), .B0(N640), .B1(N305), .Y(N944) );
  AOI22X1TF U141 ( .A0(N303), .A1(N310), .B0(N660), .B1(N302), .Y(N956) );
  AOI22X1TF U142 ( .A0(N278), .A1(N289), .B0(N682), .B1(N277), .Y(N1002) );
  AOI22X1TF U143 ( .A0(N303), .A1(N308), .B0(N662), .B1(N302), .Y(N958) );
  AOI22X1TF U144 ( .A0(N307), .A1(N306), .B0(N639), .B1(N305), .Y(N943) );
  OAI22X1TF U145 ( .A0(N642), .A1(N1640), .B0(N674), .B1(N1147), .Y(N810) );
  AOI22X1TF U146 ( .A0(N283), .A1(N289), .B0(N650), .B1(N282), .Y(N986) );
  OAI22X1TF U147 ( .A0(N641), .A1(N1640), .B0(N673), .B1(N1147), .Y(N387) );
  AOI22X1TF U148 ( .A0(N283), .A1(N293), .B0(N647), .B1(N282), .Y(N983) );
  AOI22X1TF U149 ( .A0(N280), .A1(N286), .B0(N669), .B1(N279), .Y(N997) );
  AOI22X1TF U150 ( .A0(N280), .A1(N291), .B0(N664), .B1(N279), .Y(N992) );
  AOI22X1TF U151 ( .A0(N307), .A1(N312), .B0(N642), .B1(N305), .Y(N946) );
  OAI22X1TF U152 ( .A0(N639), .A1(N1640), .B0(N671), .B1(N1147), .Y(N375) );
  AOI22X1TF U153 ( .A0(N278), .A1(N291), .B0(N680), .B1(N277), .Y(N1000) );
  AOI22X1TF U154 ( .A0(N303), .A1(N311), .B0(N659), .B1(N302), .Y(N955) );
  AOI22X1TF U155 ( .A0(N280), .A1(N293), .B0(N663), .B1(N279), .Y(N991) );
  AOI22X1TF U156 ( .A0(N298), .A1(N308), .B0(N694), .B1(N297), .Y(N974) );
  AOI22X1TF U157 ( .A0(N298), .A1(N315), .B0(N688), .B1(N297), .Y(N968) );
  AOI22X1TF U158 ( .A0(N276), .A1(N286), .B0(N701), .B1(N275), .Y(N1013) );
  NAND4XLTF U159 ( .A(N355), .B(N255), .C(N350), .D(N738), .Y(N584) );
  OAI22X1TF U160 ( .A0(N156), .A1(N620), .B0(N686), .B1(N1041), .Y(N1046) );
  AOI22X1TF U161 ( .A0(N298), .A1(N311), .B0(N691), .B1(N297), .Y(N971) );
  OAI22X1TF U162 ( .A0(N156), .A1(N608), .B0(N674), .B1(N1041), .Y(N928) );
  AOI22X1TF U163 ( .A0(N276), .A1(N291), .B0(N696), .B1(N275), .Y(N1008) );
  AOI22X1TF U164 ( .A0(N276), .A1(N289), .B0(N698), .B1(N275), .Y(N1010) );
  OAI22X1TF U165 ( .A0(N157), .A1(N607), .B0(N673), .B1(N1041), .Y(N925) );
  OAI22X1TF U166 ( .A0(N157), .A1(N6120), .B0(N678), .B1(N1041), .Y(N1021) );
  OAI22X1TF U167 ( .A0(N156), .A1(N610), .B0(N676), .B1(N1041), .Y(N934) );
  OAI22X1TF U168 ( .A0(N157), .A1(N606), .B0(N672), .B1(N1041), .Y(N922) );
  OAI22X1TF U169 ( .A0(N629), .A1(N1156), .B0(N661), .B1(N1151), .Y(N813) );
  OAI22X1TF U170 ( .A0(N625), .A1(N1156), .B0(N657), .B1(N1151), .Y(N386) );
  OAI22X1TF U171 ( .A0(N626), .A1(N1156), .B0(N658), .B1(N1151), .Y(N809) );
  OAI211X1TF U172 ( .A0(N880), .A1(N868), .B0(N871), .C0(N872), .Y(N1134) );
  NAND2BX2TF U173 ( .AN(N884), .B(N155), .Y(N1041) );
  AND3X2TF U174 ( .A(OPER3_R3[0]), .B(N371), .C(OPER3_R3[1]), .Y(N1148) );
  NAND2BX2TF U175 ( .AN(N885), .B(N155), .Y(N1044) );
  NAND4X2TF U176 ( .A(N228), .B(N239), .C(N223), .D(N371), .Y(N1146) );
  AND2X2TF U177 ( .A(\OPER1_R1[2] ), .B(N156), .Y(N174) );
  AND2X2TF U178 ( .A(N886), .B(N155), .Y(N1043) );
  AND2X2TF U179 ( .A(N355), .B(N868), .Y(N788) );
  INVX2TF U180 ( .A(N791), .Y(N126) );
  INVX1TF U181 ( .A(N842), .Y(N843) );
  OAI211XLTF U182 ( .A0(N346), .A1(N345), .B0(N558), .C0(N344), .Y(
        NEXT_STATE[2]) );
  INVX1TF U183 ( .A(N767), .Y(N769) );
  AOI22X1TF U184 ( .A0(N158), .A1(REG_A[14]), .B0(N572), .B1(REG_A[13]), .Y(
        N428) );
  NAND2XLTF U185 ( .A(REG_B[3]), .B(N590), .Y(N459) );
  AOI32X1TF U186 ( .A0(N1049), .A1(N123), .A2(N207), .B0(N268), .B1(N123), .Y(
        N269) );
  INVX2TF U187 ( .A(N1144), .Y(N130) );
  NOR2X1TF U188 ( .A(N125), .B(N582), .Y(N883) );
  NAND2XLTF U189 ( .A(N548), .B(REG_A[4]), .Y(N351) );
  INVX1TF U190 ( .A(N1050), .Y(N251) );
  INVX1TF U191 ( .A(N337), .Y(N339) );
  NAND3XLTF U192 ( .A(N861), .B(N859), .C(N208), .Y(N257) );
  INVX2TF U193 ( .A(N1172), .Y(N120) );
  INVX2TF U194 ( .A(N121), .Y(I_ADDR[0]) );
  INVX2TF U195 ( .A(N124), .Y(N125) );
  INVX2TF U196 ( .A(N791), .Y(N127) );
  INVX2TF U197 ( .A(N273), .Y(N128) );
  INVX2TF U198 ( .A(N273), .Y(N129) );
  INVX2TF U199 ( .A(N1144), .Y(N131) );
  INVX2TF U200 ( .A(N805), .Y(N132) );
  INVX2TF U201 ( .A(N805), .Y(N133) );
  INVX2TF U202 ( .A(N208), .Y(N134) );
  INVX2TF U203 ( .A(N1157), .Y(N135) );
  INVX2TF U204 ( .A(N1157), .Y(N136) );
  INVX2TF U205 ( .A(N788), .Y(N137) );
  INVX2TF U206 ( .A(N788), .Y(N138) );
  INVX2TF U207 ( .A(N130), .Y(N139) );
  INVX2TF U208 ( .A(N1137), .Y(N140) );
  INVX2TF U209 ( .A(N1137), .Y(N141) );
  INVX2TF U210 ( .A(N1134), .Y(N142) );
  INVX2TF U211 ( .A(N142), .Y(N143) );
  INVX2TF U212 ( .A(N142), .Y(N144) );
  INVX2TF U213 ( .A(N1135), .Y(N145) );
  INVX2TF U214 ( .A(N1135), .Y(N146) );
  INVX2TF U215 ( .A(N147), .Y(N148) );
  INVX2TF U216 ( .A(N147), .Y(N149) );
  INVX2TF U217 ( .A(N1043), .Y(N150) );
  INVX2TF U218 ( .A(N1043), .Y(N151) );
  INVX2TF U219 ( .A(N752), .Y(N152) );
  INVX2TF U220 ( .A(N752), .Y(N153) );
  INVX2TF U221 ( .A(N1042), .Y(N155) );
  INVX2TF U222 ( .A(N1042), .Y(N156) );
  INVX2TF U223 ( .A(N1042), .Y(N157) );
  NOR3BX1TF U224 ( .AN(N349), .B(CODE_TYPE[3]), .C(N225), .Y(N895) );
  NAND2X1TF U225 ( .A(N208), .B(N203), .Y(N349) );
  NOR2X2TF U226 ( .A(STATE[1]), .B(N230), .Y(N346) );
  AOI22X2TF U227 ( .A0(D_ADDR[8]), .A1(N129), .B0(N341), .B1(D_DATAIN[7]), .Y(
        N293) );
  OAI21X2TF U228 ( .A0(N864), .A1(N863), .B0(N862), .Y(N871) );
  NOR2X1TF U229 ( .A(CODE_TYPE[4]), .B(N358), .Y(N864) );
  AOI22X2TF U230 ( .A0(D_ADDR[6]), .A1(N128), .B0(N341), .B1(D_DATAIN[5]), .Y(
        N290) );
  AOI22X2TF U231 ( .A0(D_ADDR[4]), .A1(N128), .B0(N341), .B1(D_DATAIN[3]), .Y(
        N288) );
  AOI22X2TF U232 ( .A0(D_ADDR[1]), .A1(N129), .B0(N341), .B1(D_DATAIN[0]), .Y(
        N285) );
  AOI22X2TF U233 ( .A0(D_ADDR[3]), .A1(N129), .B0(N341), .B1(D_DATAIN[2]), .Y(
        N287) );
  AOI22X2TF U234 ( .A0(D_ADDR[5]), .A1(N129), .B0(N341), .B1(D_DATAIN[4]), .Y(
        N289) );
  AOI22X2TF U235 ( .A0(D_ADDR[7]), .A1(N129), .B0(N341), .B1(D_DATAIN[6]), .Y(
        N291) );
  AOI2BB2X2TF U236 ( .B0(D_DATAIN[7]), .B1(N296), .A0N(N412), .A1N(N295), .Y(
        N306) );
  AOI2BB2X2TF U237 ( .B0(D_DATAIN[4]), .B1(N296), .A0N(N423), .A1N(N295), .Y(
        N312) );
  AOI2BB2X2TF U238 ( .B0(D_DATAIN[5]), .B1(N296), .A0N(N420), .A1N(N295), .Y(
        N313) );
  AOI2BB2X2TF U239 ( .B0(D_DATAIN[1]), .B1(N296), .A0N(N424), .A1N(N295), .Y(
        N309) );
  AOI2BB2X2TF U240 ( .B0(D_DATAIN[2]), .B1(N296), .A0N(N421), .A1N(N295), .Y(
        N310) );
  AOI2BB2X2TF U241 ( .B0(D_DATAIN[6]), .B1(N296), .A0N(N417), .A1N(N295), .Y(
        N315) );
  AOI2BB2X2TF U242 ( .B0(D_DATAIN[3]), .B1(N296), .A0N(N418), .A1N(N295), .Y(
        N311) );
  NOR3X4TF U243 ( .A(N25), .B(N582), .C(N281), .Y(N283) );
  NOR3X4TF U244 ( .A(N125), .B(N582), .C(N304), .Y(N307) );
  NOR3X4TF U245 ( .A(N125), .B(N222), .C(N304), .Y(N303) );
  INVX2TF U246 ( .A(N24), .Y(N158) );
  INVX2TF U247 ( .A(N24), .Y(N159) );
  INVX2TF U248 ( .A(N898), .Y(N160) );
  INVX2TF U249 ( .A(N898), .Y(N161) );
  INVX2TF U250 ( .A(N899), .Y(N1620) );
  INVX2TF U251 ( .A(N899), .Y(N1630) );
  INVX2TF U252 ( .A(N1148), .Y(N1640) );
  INVX2TF U253 ( .A(N1148), .Y(N165) );
  CLKBUFX2TF U254 ( .A(N119), .Y(N245) );
  INVX2TF U255 ( .A(N738), .Y(N166) );
  NOR2X1TF U256 ( .A(N860), .B(N891), .Y(N789) );
  INVX2TF U257 ( .A(N920), .Y(N167) );
  CLKBUFX2TF U258 ( .A(N1146), .Y(N168) );
  NOR2X2TF U259 ( .A(N208), .B(N1129), .Y(N1159) );
  CLKBUFX2TF U260 ( .A(N1136), .Y(N170) );
  CLKBUFX2TF U261 ( .A(N244), .Y(N171) );
  CLKBUFX2TF U262 ( .A(N790), .Y(N244) );
  INVX2TF U263 ( .A(N839), .Y(N172) );
  NAND2X1TF U264 ( .A(N371), .B(OPER3_R3[2]), .Y(N1156) );
  NOR2X2TF U265 ( .A(N225), .B(N203), .Y(N893) );
  OAI22XLTF U266 ( .A0(N624), .A1(N172), .B0(N656), .B1(N1151), .Y(N378) );
  OAI22XLTF U267 ( .A0(N623), .A1(N1156), .B0(N655), .B1(N1151), .Y(N374) );
  OAI22XLTF U268 ( .A0(N627), .A1(N1156), .B0(N659), .B1(N1151), .Y(N382) );
  OAI22XLTF U269 ( .A0(N640), .A1(N1640), .B0(N672), .B1(N1147), .Y(N379) );
  OAI22XLTF U270 ( .A0(N645), .A1(N1640), .B0(N677), .B1(N1147), .Y(N814) );
  OAI22XLTF U271 ( .A0(N643), .A1(N1640), .B0(N675), .B1(N1147), .Y(N383) );
  NOR2X2TF U272 ( .A(CODE_TYPE[2]), .B(N579), .Y(N861) );
  INVX2TF U273 ( .A(N600), .Y(N173) );
  AOI22X2TF U274 ( .A0(D_ADDR[2]), .A1(N129), .B0(N341), .B1(D_DATAIN[1]), .Y(
        N286) );
  AOI2BB2X2TF U275 ( .B0(D_DATAIN[0]), .B1(N296), .A0N(N429), .A1N(N295), .Y(
        N308) );
  INVX2TF U276 ( .A(N174), .Y(N175) );
  INVX2TF U277 ( .A(N174), .Y(N176) );
  OAI31X4TF U278 ( .A0(N368), .A1(N348), .A2(N864), .B0(N131), .Y(N918) );
  AOI21XLTF U279 ( .A0(N1050), .A1(N346), .B0(N332), .Y(N336) );
  NOR2X2TF U280 ( .A(N207), .B(N226), .Y(N1050) );
  OAI32X4TF U281 ( .A0(N880), .A1(N857), .A2(N892), .B0(N856), .B1(N880), .Y(
        N870) );
  CLKBUFX2TF U282 ( .A(N1041), .Y(N177) );
  CLKBUFX2TF U283 ( .A(N1044), .Y(N178) );
  NOR3X4TF U284 ( .A(N25), .B(N222), .C(N281), .Y(N280) );
  CLKBUFX2TF U285 ( .A(N1149), .Y(N179) );
  CMPR32X2TF U286 ( .A(REG_A[1]), .B(REG_B[1]), .C(ADD_X_283_3_N16), .CO(
        ADD_X_283_3_N15), .S(N467) );
  CMPR32X2TF U287 ( .A(REG_A[4]), .B(REG_B[4]), .C(ADD_X_283_3_N13), .CO(
        ADD_X_283_3_N12), .S(N470) );
  CMPR32X2TF U288 ( .A(REG_A[12]), .B(REG_B[12]), .C(ADD_X_283_3_N5), .CO(
        ADD_X_283_3_N4), .S(N478) );
  CMPR32X2TF U289 ( .A(REG_A[13]), .B(REG_B[13]), .C(ADD_X_283_3_N4), .CO(
        ADD_X_283_3_N3), .S(N479) );
  ADDFHX4TF U290 ( .A(REG_A[10]), .B(REG_B[10]), .CI(ADD_X_283_3_N7), .CO(
        ADD_X_283_3_N6), .S(N476) );
  ADDFHX4TF U291 ( .A(REG_A[11]), .B(REG_B[11]), .CI(ADD_X_283_3_N6), .CO(
        ADD_X_283_3_N5), .S(N477) );
  ADDFHX2TF U292 ( .A(REG_A[3]), .B(REG_B[3]), .CI(ADD_X_283_3_N14), .CO(
        ADD_X_283_3_N13), .S(N469) );
  ADDFHX2TF U293 ( .A(REG_A[2]), .B(REG_B[2]), .CI(ADD_X_283_3_N15), .CO(
        ADD_X_283_3_N14), .S(N468) );
  ADDFHX2TF U294 ( .A(REG_A[8]), .B(REG_B[8]), .CI(ADD_X_283_3_N9), .CO(
        ADD_X_283_3_N8), .S(N474) );
  ADDFHX2TF U295 ( .A(REG_A[9]), .B(REG_B[9]), .CI(ADD_X_283_3_N8), .CO(
        ADD_X_283_3_N7), .S(N475) );
  XOR2X1TF U296 ( .A(REG_A[0]), .B(REG_B[0]), .Y(N500) );
  INVX2TF U297 ( .A(SUB_X_283_4_N1), .Y(N516) );
  CMPR32X2TF U298 ( .A(N191), .B(REG_A[12]), .C(SUB_X_283_4_N5), .CO(
        SUB_X_283_4_N4), .S(N512) );
  CMPR32X2TF U299 ( .A(N185), .B(REG_A[6]), .C(SUB_X_283_4_N11), .CO(
        SUB_X_283_4_N10), .S(N506) );
  ADDFHX4TF U300 ( .A(N189), .B(REG_A[10]), .CI(SUB_X_283_4_N7), .CO(
        SUB_X_283_4_N6), .S(N510) );
  ADDFHX4TF U301 ( .A(N190), .B(REG_A[11]), .CI(SUB_X_283_4_N6), .CO(
        SUB_X_283_4_N5), .S(N511) );
  ADDFHX4TF U302 ( .A(N194), .B(REG_A[15]), .CI(SUB_X_283_4_N2), .CO(
        SUB_X_283_4_N1), .S(N515) );
  ADDFHX2TF U303 ( .A(N193), .B(REG_A[14]), .CI(SUB_X_283_4_N3), .CO(
        SUB_X_283_4_N2), .S(N514) );
  ADDFHX4TF U304 ( .A(N187), .B(REG_A[8]), .CI(SUB_X_283_4_N9), .CO(
        SUB_X_283_4_N8), .S(N508) );
  ADDFHX4TF U305 ( .A(N188), .B(REG_A[9]), .CI(SUB_X_283_4_N8), .CO(
        SUB_X_283_4_N7), .S(N509) );
  AOI22X4TF U306 ( .A0(N514), .A1(N244), .B0(N480), .B1(N148), .Y(N405) );
  XNOR2X4TF U307 ( .A(N1168), .B(N1167), .Y(N1171) );
  AOI22X4TF U308 ( .A0(N1166), .A1(N1165), .B0(N1164), .B1(N1163), .Y(N1167)
         );
  NAND4X6TF U309 ( .A(N364), .B(N363), .C(N362), .D(N361), .Y(N1164) );
  NOR4BX4TF U310 ( .AN(N413), .B(N411), .C(N410), .D(N409), .Y(N1142) );
  AOI22X4TF U311 ( .A0(N515), .A1(N171), .B0(N481), .B1(N149), .Y(N364) );
  OAI22X1TF U312 ( .A0(N918), .A1(N1165), .B0(N919), .B1(N234), .Y(N442) );
  AOI22X2TF U313 ( .A0(N1172), .A1(N1171), .B0(N1170), .B1(N1169), .Y(N1173)
         );
  NOR3X2TF U314 ( .A(N134), .B(N358), .C(N881), .Y(N590) );
  NOR2X1TF U315 ( .A(N225), .B(N349), .Y(N366) );
  AOI221XLTF U316 ( .A0(CODE_TYPE[4]), .A1(N208), .B0(N892), .B1(N26), .C0(
        N203), .Y(N271) );
  AOI21X1TF U317 ( .A0(STATE[0]), .A1(N365), .B0(N562), .Y(N268) );
  OAI21X1TF U318 ( .A0(N893), .A1(N858), .B0(N859), .Y(N367) );
  AOI32X1TF U319 ( .A0(N893), .A1(N208), .A2(CF), .B0(N26), .B1(N258), .Y(N259) );
  AO21X1TF U320 ( .A0(N1172), .A1(N1169), .B0(N1133), .Y(N539) );
  OAI211X1TF U321 ( .A0(N749), .A1(N748), .B0(N747), .C0(N746), .Y(N1169) );
  CLKINVX4TF U322 ( .A(N1164), .Y(N1165) );
  AOI222XLTF U323 ( .A0(N737), .A1(N780), .B0(N736), .B1(N776), .C0(N766), 
        .C1(N779), .Y(N749) );
  NAND2X2TF U324 ( .A(N1162), .B(N1161), .Y(N1160) );
  NOR2X2TF U325 ( .A(CODE_TYPE[4]), .B(CODE_TYPE[3]), .Y(N859) );
  AOI31X1TF U326 ( .A0(N346), .A1(START), .A2(N207), .B0(N129), .Y(N253) );
  NAND3BX2TF U327 ( .AN(N369), .B(N1145), .C(N832), .Y(N1149) );
  NAND2X1TF U328 ( .A(N299), .B(N227), .Y(N304) );
  NAND2X1TF U329 ( .A(N227), .B(N284), .Y(N281) );
  NOR2X1TF U330 ( .A(N134), .B(CODE_TYPE[2]), .Y(N858) );
  NOR2X1TF U331 ( .A(CODE_TYPE[3]), .B(N205), .Y(N894) );
  NAND2X1TF U332 ( .A(N820), .B(N369), .Y(N372) );
  AOI21X1TF U333 ( .A0(N272), .A1(N295), .B0(N273), .Y(N299) );
  OAI22X1TF U334 ( .A0(N273), .A1(N295), .B0(N272), .B1(N274), .Y(N284) );
  NAND3X1TF U335 ( .A(N579), .B(N859), .C(N858), .Y(N272) );
  NAND2X1TF U336 ( .A(N365), .B(N1050), .Y(N274) );
  INVX2TF U337 ( .A(N252), .Y(N365) );
  NAND2X1TF U338 ( .A(N230), .B(STATE[1]), .Y(N252) );
  NOR3X4TF U339 ( .A(REG_B[2]), .B(REG_B[3]), .C(N748), .Y(N792) );
  OAI21X1TF U340 ( .A0(N562), .A1(N365), .B0(N253), .Y(N162) );
  INVX2TF U341 ( .A(N920), .Y(N1047) );
  NAND2X1TF U342 ( .A(N883), .B(N155), .Y(N920) );
  NOR2X2TF U343 ( .A(N884), .B(N304), .Y(N301) );
  NOR2BX2TF U344 ( .AN(N299), .B(N885), .Y(N298) );
  NOR2BX2TF U345 ( .AN(N284), .B(N885), .Y(N276) );
  NAND3X1TF U346 ( .A(N582), .B(N125), .C(N227), .Y(N885) );
  NOR2X2TF U347 ( .A(N884), .B(N281), .Y(N278) );
  NAND2X1TF U348 ( .A(N125), .B(N222), .Y(N884) );
  INVX2TF U349 ( .A(N274), .Y(N341) );
  INVX2TF U350 ( .A(N1170), .Y(N1143) );
  AOI211X4TF U351 ( .A0(REG_A[12]), .A1(N787), .B0(N786), .C0(N785), .Y(N1161)
         );
  AOI211X4TF U352 ( .A0(N513), .A1(N244), .B0(N764), .C0(N763), .Y(N1162) );
  NOR2X1TF U353 ( .A(N205), .B(N229), .Y(N855) );
  NAND3X1TF U354 ( .A(CODE_TYPE[2]), .B(N134), .C(N203), .Y(N891) );
  AO22X1TF U355 ( .A0(N256), .A1(N482), .B0(N516), .B1(N171), .Y(N585) );
  NAND2X1TF U356 ( .A(N230), .B(N1050), .Y(N344) );
  AOI222XLTF U357 ( .A0(N267), .A1(N328), .B0(I_ADDR[8]), .B1(N331), .C0(
        D_ADDR[8]), .C1(N330), .Y(N873) );
  NOR2X1TF U358 ( .A(N327), .B(N233), .Y(N334) );
  NAND2X1TF U359 ( .A(N855), .B(N262), .Y(N265) );
  NAND2X1TF U360 ( .A(N329), .B(I_ADDR[7]), .Y(N327) );
  INVX2TF U361 ( .A(N1054), .Y(N1053) );
  NAND2X2TF U362 ( .A(N1050), .B(N1049), .Y(N1054) );
  INVX2TF U363 ( .A(N917), .Y(N916) );
  NAND2X2TF U364 ( .A(N906), .B(N1049), .Y(N917) );
  INVX2TF U365 ( .A(N345), .Y(N906) );
  INVX2TF U366 ( .A(N301), .Y(N300) );
  INVX2TF U367 ( .A(N303), .Y(N302) );
  INVX2TF U368 ( .A(N298), .Y(N297) );
  INVX2TF U369 ( .A(N307), .Y(N305) );
  INVX2TF U370 ( .A(N272), .Y(N296) );
  INVX2TF U371 ( .A(N314), .Y(N316) );
  INVX2TF U372 ( .A(N276), .Y(N275) );
  INVX2TF U373 ( .A(N283), .Y(N282) );
  INVX2TF U374 ( .A(N278), .Y(N277) );
  INVX2TF U375 ( .A(N280), .Y(N279) );
  INVX2TF U376 ( .A(N292), .Y(N294) );
  AND2X2TF U377 ( .A(STATE[1]), .B(N564), .Y(N1049) );
  NAND2X1TF U378 ( .A(N346), .B(N1050), .Y(N340) );
  NAND2X1TF U379 ( .A(N173), .B(REG_A[15]), .Y(N801) );
  NAND2X1TF U380 ( .A(N173), .B(REG_A[5]), .Y(N427) );
  INVX2TF U381 ( .A(N789), .Y(N738) );
  NAND2X1TF U382 ( .A(N152), .B(REG_A[5]), .Y(N5850) );
  NAND2X1TF U383 ( .A(N152), .B(REG_A[8]), .Y(N5000) );
  AOI21X1TF U384 ( .A0(N572), .A1(REG_A[2]), .B0(N394), .Y(N441) );
  NAND2X1TF U385 ( .A(N572), .B(REG_A[6]), .Y(N491) );
  NAND2X1TF U386 ( .A(N572), .B(REG_A[0]), .Y(N775) );
  AOI211X1TF U387 ( .A0(N894), .A1(N366), .B0(N890), .C0(N126), .Y(N355) );
  NOR2X1TF U388 ( .A(N881), .B(N891), .Y(N890) );
  NOR2X1TF U389 ( .A(N249), .B(N171), .Y(N255) );
  AOI21X1TF U390 ( .A0(N343), .A1(N342), .B0(N341), .Y(N558) );
  OAI21X1TF U391 ( .A0(N340), .A1(N339), .B0(N338), .Y(N342) );
  OAI31X1TF U392 ( .A0(N208), .A1(N882), .A2(N881), .B0(N128), .Y(N333) );
  NOR2X1TF U393 ( .A(IO_STATUS[0]), .B(IO_STATUS[1]), .Y(N343) );
  OAI21X1TF U394 ( .A0(N647), .A1(N920), .B0(N905), .Y(N462) );
  AOI211X1TF U395 ( .A0(N174), .A1(IO_OFFSET[7]), .B0(N904), .C0(N903), .Y(
        N905) );
  OAI22X1TF U396 ( .A0(N695), .A1(N178), .B0(N663), .B1(N151), .Y(N903) );
  OAI22X1TF U397 ( .A0(N157), .A1(N613), .B0(N679), .B1(N177), .Y(N904) );
  OAI21X1TF U398 ( .A0(N651), .A1(N920), .B0(N889), .Y(N458) );
  AOI211X1TF U399 ( .A0(N174), .A1(IO_OFFSET[3]), .B0(N888), .C0(N887), .Y(
        N889) );
  OAI22X1TF U400 ( .A0(N699), .A1(N178), .B0(N667), .B1(N151), .Y(N887) );
  OAI22X1TF U401 ( .A0(N156), .A1(N617), .B0(N683), .B1(N177), .Y(N888) );
  AOI211X1TF U402 ( .A0(N1047), .A1(IO_DATAOUTB[0]), .B0(N1046), .C0(N1045), 
        .Y(N1048) );
  OAI22X1TF U403 ( .A0(N697), .A1(N178), .B0(N665), .B1(N150), .Y(N1029) );
  OAI22X1TF U404 ( .A0(N157), .A1(N615), .B0(N681), .B1(N177), .Y(N1030) );
  OAI22X1TF U405 ( .A0(N687), .A1(N178), .B0(N655), .B1(N150), .Y(N1023) );
  OAI22X1TF U406 ( .A0(N156), .A1(N605), .B0(N671), .B1(N177), .Y(N1024) );
  OAI22X1TF U407 ( .A0(N701), .A1(N178), .B0(N669), .B1(N151), .Y(N1038) );
  OAI22X1TF U408 ( .A0(N157), .A1(N619), .B0(N685), .B1(N177), .Y(N1039) );
  OAI22X1TF U409 ( .A0(N693), .A1(N178), .B0(N661), .B1(N151), .Y(N1017) );
  OAI22X1TF U410 ( .A0(N156), .A1(N611), .B0(N677), .B1(N177), .Y(N1018) );
  OAI22X1TF U411 ( .A0(N700), .A1(N178), .B0(N668), .B1(N151), .Y(N1035) );
  OAI22X1TF U412 ( .A0(N157), .A1(N618), .B0(N684), .B1(N177), .Y(N1036) );
  OAI22X1TF U413 ( .A0(N691), .A1(N178), .B0(N659), .B1(N151), .Y(N930) );
  OAI22X1TF U414 ( .A0(N156), .A1(N609), .B0(N675), .B1(N177), .Y(N931) );
  OAI22X1TF U415 ( .A0(N696), .A1(N178), .B0(N664), .B1(N151), .Y(N1026) );
  OAI22X1TF U416 ( .A0(N157), .A1(N614), .B0(N680), .B1(N177), .Y(N1027) );
  OAI22X1TF U417 ( .A0(N698), .A1(N178), .B0(N666), .B1(N151), .Y(N1032) );
  OAI22X1TF U418 ( .A0(N156), .A1(N616), .B0(N682), .B1(N177), .Y(N1033) );
  INVX2TF U419 ( .A(N918), .Y(N919) );
  OAI21X1TF U420 ( .A0(N635), .A1(N172), .B0(N851), .Y(N456) );
  NOR3X1TF U421 ( .A(N850), .B(N849), .C(N848), .Y(N851) );
  OAI22X1TF U422 ( .A0(N667), .A1(N247), .B0(N182), .B1(N1149), .Y(N848) );
  OAI22X1TF U423 ( .A0(N651), .A1(N165), .B0(N683), .B1(N246), .Y(N849) );
  OAI22X1TF U424 ( .A0(N699), .A1(N168), .B0(N431), .B1(N1145), .Y(N850) );
  NOR3X1TF U425 ( .A(N846), .B(N845), .C(N844), .Y(N847) );
  OAI22X1TF U426 ( .A0(N663), .A1(N247), .B0(N186), .B1(N1149), .Y(N844) );
  OAI22X1TF U427 ( .A0(N647), .A1(N1640), .B0(N679), .B1(N246), .Y(N845) );
  OAI22X1TF U428 ( .A0(N432), .A1(N843), .B0(N695), .B1(N1146), .Y(N846) );
  OAI21X1TF U429 ( .A0(N190), .A1(N1149), .B0(N385), .Y(N445) );
  NOR3X1TF U430 ( .A(N384), .B(N383), .C(N382), .Y(N385) );
  OAI22X1TF U431 ( .A0(N691), .A1(N1146), .B0(N431), .B1(N832), .Y(N384) );
  OAI21X1TF U432 ( .A0(N194), .A1(N179), .B0(N377), .Y(N443) );
  NOR3X1TF U433 ( .A(N376), .B(N375), .C(N374), .Y(N377) );
  OAI22X1TF U434 ( .A0(N687), .A1(N1146), .B0(N432), .B1(N832), .Y(N376) );
  OAI21X1TF U435 ( .A0(N191), .A1(N179), .B0(N812), .Y(N449) );
  NOR3X1TF U436 ( .A(N811), .B(N810), .C(N809), .Y(N812) );
  OAI22X1TF U437 ( .A0(N690), .A1(N1146), .B0(N416), .B1(N832), .Y(N811) );
  OAI21X1TF U438 ( .A0(N187), .A1(N179), .B0(N836), .Y(N453) );
  NOR3X1TF U439 ( .A(N835), .B(N834), .C(N833), .Y(N836) );
  OAI22X1TF U440 ( .A0(N630), .A1(N172), .B0(N662), .B1(N247), .Y(N833) );
  OAI22X1TF U441 ( .A0(N646), .A1(N165), .B0(N678), .B1(N246), .Y(N834) );
  OAI22X1TF U442 ( .A0(N694), .A1(N1146), .B0(N228), .B1(N832), .Y(N835) );
  OAI21X1TF U443 ( .A0(N192), .A1(N179), .B0(N389), .Y(N446) );
  NOR3X1TF U444 ( .A(N388), .B(N387), .C(N386), .Y(N389) );
  OAI22X1TF U445 ( .A0(N689), .A1(N1146), .B0(N415), .B1(N832), .Y(N388) );
  OAI21X1TF U446 ( .A0(N189), .A1(N179), .B0(N393), .Y(N447) );
  NOR3X1TF U447 ( .A(N392), .B(N391), .C(N390), .Y(N393) );
  OAI22X1TF U448 ( .A0(N628), .A1(N172), .B0(N660), .B1(N247), .Y(N390) );
  OAI22X1TF U449 ( .A0(N644), .A1(N165), .B0(N676), .B1(N246), .Y(N391) );
  OAI22X1TF U450 ( .A0(N692), .A1(N168), .B0(N239), .B1(N832), .Y(N392) );
  OAI21X1TF U451 ( .A0(N188), .A1(N179), .B0(N816), .Y(N450) );
  NOR3X1TF U452 ( .A(N815), .B(N814), .C(N813), .Y(N816) );
  OAI22X1TF U453 ( .A0(N693), .A1(N168), .B0(N223), .B1(N832), .Y(N815) );
  OAI21X1TF U454 ( .A0(N193), .A1(N179), .B0(N381), .Y(N444) );
  NOR3X1TF U455 ( .A(N380), .B(N379), .C(N378), .Y(N381) );
  OAI22X1TF U456 ( .A0(N688), .A1(N168), .B0(N414), .B1(N832), .Y(N380) );
  NOR3X1TF U457 ( .A(N1094), .B(N1093), .C(N1092), .Y(N1095) );
  OAI22X1TF U458 ( .A0(N668), .A1(N247), .B0(N181), .B1(N1149), .Y(N1092) );
  OAI22X1TF U459 ( .A0(N652), .A1(N1640), .B0(N684), .B1(N246), .Y(N1093) );
  OAI22X1TF U460 ( .A0(N700), .A1(N1146), .B0(N239), .B1(N1145), .Y(N1094) );
  NOR3X1TF U461 ( .A(N1127), .B(N1126), .C(N1125), .Y(N1128) );
  OAI22X1TF U462 ( .A0(N669), .A1(N247), .B0(N1124), .B1(N1149), .Y(N1125) );
  OAI22X1TF U463 ( .A0(N653), .A1(N165), .B0(N685), .B1(N246), .Y(N1126) );
  OAI22X1TF U464 ( .A0(N701), .A1(N1146), .B0(N223), .B1(N1145), .Y(N1127) );
  NOR3X1TF U465 ( .A(N1154), .B(N1153), .C(N1152), .Y(N1155) );
  OAI22X1TF U466 ( .A0(N670), .A1(N247), .B0(N1150), .B1(N1149), .Y(N1152) );
  OAI22X1TF U467 ( .A0(N654), .A1(N165), .B0(N686), .B1(N246), .Y(N1153) );
  OAI22X1TF U468 ( .A0(N702), .A1(N1146), .B0(N228), .B1(N1145), .Y(N1154) );
  OAI211X1TF U469 ( .A0(N697), .A1(N168), .B0(N841), .C0(N840), .Y(N454) );
  AOI211X1TF U470 ( .A0(N839), .A1(IO_OFFSET[5]), .B0(N838), .C0(N837), .Y(
        N841) );
  OAI22X1TF U471 ( .A0(N665), .A1(N247), .B0(N184), .B1(N1149), .Y(N837) );
  OAI22X1TF U472 ( .A0(N649), .A1(N165), .B0(N681), .B1(N246), .Y(N838) );
  OAI211X1TF U473 ( .A0(N696), .A1(N168), .B0(N831), .C0(N830), .Y(N452) );
  AOI211X1TF U474 ( .A0(N839), .A1(IO_OFFSET[6]), .B0(N829), .C0(N828), .Y(
        N831) );
  OAI22X1TF U475 ( .A0(N664), .A1(N247), .B0(N185), .B1(N1149), .Y(N828) );
  OAI22X1TF U476 ( .A0(N648), .A1(N165), .B0(N680), .B1(N246), .Y(N829) );
  OAI211X1TF U477 ( .A0(N698), .A1(N168), .B0(N827), .C0(N826), .Y(N451) );
  NOR2X1TF U478 ( .A(N820), .B(N880), .Y(N842) );
  AOI211X1TF U479 ( .A0(N839), .A1(IO_OFFSET[4]), .B0(N819), .C0(N818), .Y(
        N827) );
  OAI22X1TF U480 ( .A0(N666), .A1(N247), .B0(N183), .B1(N1149), .Y(N818) );
  NAND2X2TF U481 ( .A(N368), .B(N862), .Y(N832) );
  NOR2X1TF U482 ( .A(OPER3_R3[0]), .B(N372), .Y(N373) );
  OAI22X1TF U483 ( .A0(N650), .A1(N165), .B0(N682), .B1(N246), .Y(N819) );
  NOR2X1TF U484 ( .A(OPER3_R3[1]), .B(N372), .Y(N370) );
  INVX2TF U485 ( .A(N1156), .Y(N839) );
  INVX2TF U486 ( .A(N372), .Y(N371) );
  AOI211X1TF U487 ( .A0(N229), .A1(N891), .B0(N880), .C0(CODE_TYPE[4]), .Y(
        N369) );
  AOI211X1TF U488 ( .A0(CODE_TYPE[4]), .A1(N366), .B0(N855), .C0(N853), .Y(
        N820) );
  OAI21X1TF U489 ( .A0(N651), .A1(N899), .B0(N879), .Y(N457) );
  AOI211X1TF U490 ( .A0(IO_CONTROL[3]), .A1(N898), .B0(N878), .C0(N877), .Y(
        N879) );
  OAI21X1TF U491 ( .A0(N677), .A1(N160), .B0(N1087), .Y(N5160) );
  AOI211X1TF U492 ( .A0(IO_DATAOUTB[9]), .A1(N1620), .B0(N1086), .C0(N1085), 
        .Y(N1087) );
  OAI21X1TF U493 ( .A0(N678), .A1(N160), .B0(N1066), .Y(N5070) );
  AOI211X1TF U494 ( .A0(IO_DATAOUTB[8]), .A1(N1620), .B0(N1065), .C0(N1064), 
        .Y(N1066) );
  OAI21X1TF U495 ( .A0(N675), .A1(N160), .B0(N1117), .Y(N531) );
  AOI211X1TF U496 ( .A0(IO_DATAOUTB[11]), .A1(N1620), .B0(N1116), .C0(N1115), 
        .Y(N1117) );
  OAI21X1TF U497 ( .A0(N676), .A1(N160), .B0(N1106), .Y(N525) );
  AOI211X1TF U498 ( .A0(IO_DATAOUTB[10]), .A1(N1620), .B0(N1105), .C0(N1104), 
        .Y(N1106) );
  OAI21X1TF U499 ( .A0(N673), .A1(N160), .B0(N1112), .Y(N528) );
  AOI211X1TF U500 ( .A0(N240), .A1(N1620), .B0(N1111), .C0(N1110), .Y(N1112)
         );
  OAI21X1TF U501 ( .A0(N685), .A1(N160), .B0(N912), .Y(N465) );
  AOI211X1TF U502 ( .A0(IO_DATAOUTB[1]), .A1(N1620), .B0(N911), .C0(N910), .Y(
        N912) );
  OAI21X1TF U503 ( .A0(N681), .A1(N160), .B0(N1060), .Y(N5040) );
  AOI211X1TF U504 ( .A0(IO_DATAOUTB[5]), .A1(N1620), .B0(N1059), .C0(N1058), 
        .Y(N1060) );
  OAI21X1TF U505 ( .A0(N672), .A1(N160), .B0(N1123), .Y(N534) );
  AOI211X1TF U506 ( .A0(N241), .A1(N1620), .B0(N1122), .C0(N1121), .Y(N1123)
         );
  OAI21X1TF U507 ( .A0(N682), .A1(N161), .B0(N1080), .Y(N5130) );
  AOI211X1TF U508 ( .A0(IO_DATAOUTB[4]), .A1(N1630), .B0(N1079), .C0(N1078), 
        .Y(N1080) );
  OAI21X1TF U509 ( .A0(N679), .A1(N161), .B0(N902), .Y(N461) );
  AOI211X1TF U510 ( .A0(IO_DATAOUTB[7]), .A1(N1630), .B0(N901), .C0(N900), .Y(
        N902) );
  AOI211X1TF U511 ( .A0(IO_DATAOUTB[6]), .A1(N1630), .B0(N1072), .C0(N1071), 
        .Y(N1073) );
  OAI21X1TF U512 ( .A0(N671), .A1(N161), .B0(N11400), .Y(N540) );
  AOI211X1TF U513 ( .A0(N242), .A1(N1630), .B0(N1139), .C0(N1138), .Y(N11400)
         );
  OAI21X1TF U514 ( .A0(N674), .A1(N161), .B0(N1101), .Y(N522) );
  AOI211X1TF U515 ( .A0(IO_DATAOUTB[12]), .A1(N1630), .B0(N1100), .C0(N1099), 
        .Y(N1101) );
  OAI21X1TF U516 ( .A0(N684), .A1(N161), .B0(N915), .Y(N4660) );
  AOI211X1TF U517 ( .A0(IO_DATAOUTB[2]), .A1(N1630), .B0(N914), .C0(N913), .Y(
        N915) );
  OAI21X1TF U518 ( .A0(N686), .A1(N161), .B0(N909), .Y(N464) );
  AOI211X1TF U519 ( .A0(IO_DATAOUTB[0]), .A1(N1630), .B0(N908), .C0(N907), .Y(
        N909) );
  AOI31X4TF U520 ( .A0(N876), .A1(N415), .A2(N414), .B0(N875), .Y(N1136) );
  NOR2X1TF U521 ( .A(N872), .B(N885), .Y(N875) );
  NOR2X1TF U522 ( .A(N871), .B(N238), .Y(N876) );
  NOR2X1TF U523 ( .A(N415), .B(N871), .Y(N867) );
  NOR2X1TF U524 ( .A(N125), .B(N222), .Y(N886) );
  AOI22X1TF U525 ( .A0(N883), .A1(N870), .B0(N865), .B1(N237), .Y(N899) );
  NOR2X1TF U526 ( .A(N416), .B(N871), .Y(N865) );
  INVX2TF U527 ( .A(N870), .Y(N872) );
  AOI211X1TF U528 ( .A0(N855), .A1(N854), .B0(N853), .C0(N852), .Y(N856) );
  NOR2X1TF U529 ( .A(N229), .B(N882), .Y(N853) );
  INVX2TF U530 ( .A(N861), .Y(N882) );
  INVX2TF U531 ( .A(N871), .Y(N869) );
  INVX2TF U532 ( .A(N880), .Y(N862) );
  NAND2X2TF U533 ( .A(N906), .B(N365), .Y(N880) );
  AOI21X1TF U534 ( .A0(N347), .A1(N857), .B0(N892), .Y(N368) );
  AOI21X1TF U535 ( .A0(D_ADDR[1]), .A1(N330), .B0(N266), .Y(N874) );
  AOI211X1TF U536 ( .A0(N330), .A1(D_ADDR[6]), .B0(N326), .C0(N325), .Y(N821)
         );
  AOI211X1TF U537 ( .A0(N324), .A1(N232), .B0(N329), .C0(N323), .Y(N325) );
  NOR2X1TF U538 ( .A(N232), .B(N322), .Y(N326) );
  AOI211X1TF U539 ( .A0(N330), .A1(D_ADDR[4]), .B0(N320), .C0(N319), .Y(N823)
         );
  AOI211X1TF U540 ( .A0(N318), .A1(N231), .B0(N321), .C0(N323), .Y(N319) );
  NOR2X1TF U541 ( .A(N231), .B(N322), .Y(N320) );
  INVX2TF U542 ( .A(N322), .Y(N331) );
  OAI211X1TF U543 ( .A0(N334), .A1(N273), .B0(N264), .C0(N263), .Y(N322) );
  INVX2TF U544 ( .A(N330), .Y(N263) );
  NOR2X2TF U545 ( .A(N273), .B(N265), .Y(N330) );
  INVX2TF U546 ( .A(N323), .Y(N328) );
  OAI211X1TF U547 ( .A0(CF), .A1(N261), .B0(N260), .C0(N259), .Y(N262) );
  AOI32X1TF U548 ( .A0(N579), .A1(ZF), .A2(N225), .B0(N861), .B1(N235), .Y(
        N260) );
  NOR2X1TF U549 ( .A(N324), .B(N232), .Y(N329) );
  NOR2X1TF U550 ( .A(N318), .B(N231), .Y(N321) );
  AOI22X1TF U551 ( .A0(N123), .A1(N605), .B0(N613), .B1(N121), .Y(D_DATAOUT[7]) );
  AOI22X1TF U552 ( .A0(N123), .A1(N606), .B0(N614), .B1(N121), .Y(D_DATAOUT[6]) );
  AOI22X1TF U553 ( .A0(N123), .A1(N607), .B0(N615), .B1(N121), .Y(D_DATAOUT[5]) );
  AOI22X1TF U554 ( .A0(N123), .A1(N608), .B0(N616), .B1(N121), .Y(D_DATAOUT[4]) );
  AOI22X1TF U555 ( .A0(N123), .A1(N609), .B0(N617), .B1(N121), .Y(D_DATAOUT[3]) );
  AOI22X1TF U556 ( .A0(I_ADDR[0]), .A1(N610), .B0(N618), .B1(N121), .Y(
        D_DATAOUT[2]) );
  AOI22X1TF U557 ( .A0(I_ADDR[0]), .A1(N611), .B0(N619), .B1(N121), .Y(
        D_DATAOUT[1]) );
  AOI22X1TF U558 ( .A0(I_ADDR[0]), .A1(N6120), .B0(N620), .B1(N121), .Y(
        D_DATAOUT[0]) );
  AOI22X1TF U559 ( .A0(N1053), .A1(N1051), .B0(N205), .B1(N1054), .Y(N492) );
  AOI22X1TF U560 ( .A0(N1053), .A1(N1052), .B0(N579), .B1(N1054), .Y(N496) );
  AOI22X1TF U561 ( .A0(N916), .A1(N1051), .B0(N432), .B1(N917), .Y(N463) );
  INVX2TF U562 ( .A(I_DATAIN[7]), .Y(N1051) );
  AOI22X1TF U563 ( .A0(N916), .A1(N1052), .B0(N431), .B1(N917), .Y(N4700) );
  INVX2TF U564 ( .A(I_DATAIN[3]), .Y(N1052) );
  OAI211X1TF U565 ( .A0(N251), .A1(N230), .B0(N338), .C0(N335), .Y(N114) );
  INVX2TF U566 ( .A(N332), .Y(N338) );
  NOR3X1TF U567 ( .A(STATE[0]), .B(N562), .C(N252), .Y(N332) );
  AOI22X1TF U568 ( .A0(N301), .A1(N306), .B0(N671), .B1(N300), .Y(N959) );
  AOI22X1TF U569 ( .A0(N298), .A1(N306), .B0(N687), .B1(N297), .Y(N967) );
  AOI22X1TF U570 ( .A0(N298), .A1(N309), .B0(N693), .B1(N297), .Y(N973) );
  AOI22X1TF U571 ( .A0(N301), .A1(N309), .B0(N677), .B1(N300), .Y(N965) );
  AOI22X1TF U572 ( .A0(N298), .A1(N312), .B0(N690), .B1(N297), .Y(N970) );
  AOI22X1TF U573 ( .A0(N298), .A1(N310), .B0(N692), .B1(N297), .Y(N972) );
  AOI22X1TF U574 ( .A0(N298), .A1(N313), .B0(N689), .B1(N297), .Y(N969) );
  AOI22X1TF U575 ( .A0(N303), .A1(N315), .B0(N656), .B1(N302), .Y(N952) );
  AOI22X1TF U576 ( .A0(N303), .A1(N313), .B0(N657), .B1(N302), .Y(N953) );
  AOI22X1TF U577 ( .A0(N301), .A1(N313), .B0(N673), .B1(N300), .Y(N961) );
  AOI22X1TF U578 ( .A0(N301), .A1(N312), .B0(N674), .B1(N300), .Y(N962) );
  AOI22X1TF U579 ( .A0(N301), .A1(N310), .B0(N676), .B1(N300), .Y(N964) );
  AOI22X1TF U580 ( .A0(N307), .A1(N311), .B0(N643), .B1(N305), .Y(N947) );
  AOI22X1TF U581 ( .A0(N303), .A1(N312), .B0(N658), .B1(N302), .Y(N954) );
  AOI22X1TF U582 ( .A0(N307), .A1(N309), .B0(N645), .B1(N305), .Y(N949) );
  AOI22X1TF U583 ( .A0(N307), .A1(N310), .B0(N644), .B1(N305), .Y(N948) );
  AOI22X1TF U584 ( .A0(N316), .A1(N306), .B0(N623), .B1(N314), .Y(N1015) );
  AOI22X1TF U585 ( .A0(N316), .A1(N312), .B0(N626), .B1(N314), .Y(N938) );
  AOI22X1TF U586 ( .A0(N316), .A1(N308), .B0(N630), .B1(N314), .Y(N942) );
  AOI22X1TF U587 ( .A0(N316), .A1(N313), .B0(N625), .B1(N314), .Y(N937) );
  AOI22X1TF U588 ( .A0(N316), .A1(N309), .B0(N629), .B1(N314), .Y(N941) );
  AOI22X1TF U589 ( .A0(N316), .A1(N310), .B0(N628), .B1(N314), .Y(N940) );
  AOI22X1TF U590 ( .A0(N316), .A1(N315), .B0(N624), .B1(N314), .Y(N936) );
  AOI22X1TF U591 ( .A0(N316), .A1(N311), .B0(N627), .B1(N314), .Y(N939) );
  NAND4X2TF U592 ( .A(N25), .B(N582), .C(\OPER1_R1[2] ), .D(N299), .Y(N314) );
  AOI22X1TF U593 ( .A0(N278), .A1(N293), .B0(N679), .B1(N277), .Y(N999) );
  AOI22X1TF U594 ( .A0(N276), .A1(N293), .B0(N695), .B1(N275), .Y(N1007) );
  AOI22X1TF U595 ( .A0(N278), .A1(N285), .B0(N686), .B1(N277), .Y(N1006) );
  AOI22X1TF U596 ( .A0(N276), .A1(N290), .B0(N697), .B1(N275), .Y(N1009) );
  AOI22X1TF U597 ( .A0(N283), .A1(N291), .B0(N648), .B1(N282), .Y(N984) );
  AOI22X1TF U598 ( .A0(N276), .A1(N287), .B0(N700), .B1(N275), .Y(N1012) );
  AOI22X1TF U599 ( .A0(N276), .A1(N285), .B0(N702), .B1(N275), .Y(N1014) );
  AOI22X1TF U600 ( .A0(N276), .A1(N288), .B0(N699), .B1(N275), .Y(N1011) );
  AOI22X1TF U601 ( .A0(N283), .A1(N290), .B0(N649), .B1(N282), .Y(N985) );
  AOI22X1TF U602 ( .A0(N278), .A1(N287), .B0(N684), .B1(N277), .Y(N1004) );
  AOI22X1TF U603 ( .A0(N280), .A1(N287), .B0(N668), .B1(N279), .Y(N996) );
  AOI22X1TF U604 ( .A0(N278), .A1(N290), .B0(N681), .B1(N277), .Y(N1001) );
  AOI22X1TF U605 ( .A0(N278), .A1(N288), .B0(N683), .B1(N277), .Y(N1003) );
  AOI22X1TF U606 ( .A0(N280), .A1(N285), .B0(N670), .B1(N279), .Y(N998) );
  AOI22X1TF U607 ( .A0(N283), .A1(N288), .B0(N651), .B1(N282), .Y(N987) );
  AOI22X1TF U608 ( .A0(N280), .A1(N289), .B0(N666), .B1(N279), .Y(N994) );
  AOI22X1TF U609 ( .A0(N294), .A1(N293), .B0(N631), .B1(N292), .Y(N975) );
  AOI22X1TF U610 ( .A0(N294), .A1(N289), .B0(N634), .B1(N292), .Y(N978) );
  AOI22X1TF U611 ( .A0(N294), .A1(N290), .B0(N633), .B1(N292), .Y(N977) );
  AOI22X1TF U612 ( .A0(N294), .A1(N286), .B0(N637), .B1(N292), .Y(N981) );
  AOI22X1TF U613 ( .A0(N294), .A1(N285), .B0(N638), .B1(N292), .Y(N982) );
  AOI22X1TF U614 ( .A0(N294), .A1(N287), .B0(N636), .B1(N292), .Y(N980) );
  AOI22X1TF U615 ( .A0(N294), .A1(N291), .B0(N632), .B1(N292), .Y(N976) );
  AOI22X1TF U616 ( .A0(N294), .A1(N288), .B0(N635), .B1(N292), .Y(N979) );
  NAND4X2TF U617 ( .A(N582), .B(N25), .C(\OPER1_R1[2] ), .D(N284), .Y(N292) );
  OAI31X4TF U618 ( .A0(N895), .A1(N271), .A2(N270), .B0(N272), .Y(N295) );
  OAI22X1TF U619 ( .A0(N893), .A1(N860), .B0(N892), .B1(N349), .Y(N270) );
  OAI211X1TF U620 ( .A0(N1161), .A1(N1143), .B0(N1103), .C0(N1102), .Y(N524)
         );
  AOI22X1TF U621 ( .A0(IO_DATAINA[12]), .A1(N169), .B0(N1172), .B1(N1118), .Y(
        N1102) );
  OAI211X1TF U622 ( .A0(N1132), .A1(N1141), .B0(N1098), .C0(N1097), .Y(N521)
         );
  AOI22X1TF U623 ( .A0(IO_DATAINB[2]), .A1(N135), .B0(D_ADDR[3]), .B1(N139), 
        .Y(N1098) );
  OAI21X1TF U624 ( .A0(N1162), .A1(N1143), .B0(N1114), .Y(N530) );
  AOI21X1TF U625 ( .A0(N169), .A1(IO_DATAINA[13]), .B0(N1113), .Y(N1114) );
  OAI22X1TF U626 ( .A0(N1161), .A1(N1141), .B0(N131), .B1(N420), .Y(N1113) );
  OAI211X1TF U627 ( .A0(N1109), .A1(N120), .B0(N1108), .C0(N1107), .Y(N527) );
  AOI22X1TF U628 ( .A0(IO_DATAINA[10]), .A1(N1159), .B0(N1170), .B1(N1163), 
        .Y(N1107) );
  OAI211X1TF U629 ( .A0(N1096), .A1(N120), .B0(N897), .C0(N896), .Y(N460) );
  AOI22X1TF U630 ( .A0(IO_DATAINA[3]), .A1(N1159), .B0(N1170), .B1(N1081), .Y(
        N896) );
  AOI22X1TF U631 ( .A0(IO_DATAINB[3]), .A1(N135), .B0(D_ADDR[4]), .B1(N139), 
        .Y(N897) );
  OAI211X1TF U632 ( .A0(N5110), .A1(N773), .B0(N5080), .C0(N5050), .Y(N5140)
         );
  AOI22X1TF U633 ( .A0(REG_B[2]), .A1(N5020), .B0(REG_A[2]), .B1(N5010), .Y(
        N5050) );
  OAI21X1TF U634 ( .A0(REG_B[2]), .A1(N224), .B0(N592), .Y(N5010) );
  AOI22X1TF U635 ( .A0(N796), .A1(N711), .B0(N502), .B1(N244), .Y(N5080) );
  INVX2TF U636 ( .A(N490), .Y(N5110) );
  OAI211X1TF U637 ( .A0(N209), .A1(N752), .B0(N570), .C0(N565), .Y(N490) );
  OAI22X1TF U638 ( .A0(N489), .A1(N459), .B0(N441), .B1(N805), .Y(N517) );
  OAI211X1TF U639 ( .A0(N1109), .A1(N1143), .B0(N1091), .C0(N1090), .Y(N518)
         );
  AOI22X1TF U640 ( .A0(IO_DATAINA[9]), .A1(N169), .B0(N1172), .B1(N1089), .Y(
        N1090) );
  INVX2TF U641 ( .A(N1088), .Y(N1109) );
  OAI211X1TF U642 ( .A0(N188), .A1(N561), .B0(N560), .C0(N559), .Y(N1088) );
  OAI31X1TF U643 ( .A0(N182), .A1(N782), .A2(N555), .B0(N554), .Y(N556) );
  AOI22X1TF U644 ( .A0(N798), .A1(N726), .B0(N796), .B1(N725), .Y(N554) );
  OAI211X1TF U645 ( .A0(N1166), .A1(N120), .B0(N1120), .C0(N1119), .Y(N533) );
  AOI22X1TF U646 ( .A0(IO_DATAINA[11]), .A1(N1159), .B0(N1170), .B1(N1118), 
        .Y(N1119) );
  OAI211X1TF U647 ( .A0(N190), .A1(N547), .B0(N546), .C0(N544), .Y(N1118) );
  OAI21X1TF U648 ( .A0(N801), .A1(N532), .B0(N529), .Y(N535) );
  AOI22X1TF U649 ( .A0(N526), .A1(N797), .B0(N798), .B1(N804), .Y(N529) );
  INVX2TF U650 ( .A(N576), .Y(N526) );
  OAI22X1TF U651 ( .A0(N523), .A1(N220), .B0(N591), .B1(N773), .Y(N538) );
  OAI211X1TF U652 ( .A0(N1070), .A1(N120), .B0(N1069), .C0(N1068), .Y(N5090)
         );
  AOI22X1TF U653 ( .A0(IO_DATAINA[8]), .A1(N1159), .B0(N1170), .B1(N1089), .Y(
        N1068) );
  OAI211X1TF U654 ( .A0(N187), .A1(N583), .B0(N581), .C0(N580), .Y(N1089) );
  OAI21X1TF U655 ( .A0(N576), .A1(N775), .B0(N575), .Y(N577) );
  AOI22X1TF U656 ( .A0(N798), .A1(N781), .B0(N796), .B1(N766), .Y(N575) );
  OAI22X1TF U657 ( .A0(N569), .A1(N215), .B0(N622), .B1(N773), .Y(N578) );
  INVX2TF U658 ( .A(N1067), .Y(N1070) );
  OAI211X1TF U659 ( .A0(N1132), .A1(N1143), .B0(N1131), .C0(N1130), .Y(N1133)
         );
  AOI22X1TF U660 ( .A0(N1159), .A1(IO_DATAINA[1]), .B0(N1158), .B1(
        IO_STATUS[1]), .Y(N1130) );
  AOI22X1TF U661 ( .A0(IO_DATAINB[1]), .A1(N135), .B0(D_ADDR[2]), .B1(N139), 
        .Y(N1131) );
  AOI211X1TF U662 ( .A0(REG_B[1]), .A1(N440), .B0(N439), .C0(N438), .Y(N1132)
         );
  OAI211X1TF U663 ( .A0(N437), .A1(N748), .B0(N436), .C0(N435), .Y(N438) );
  OAI211X1TF U664 ( .A0(N209), .A1(N119), .B0(N433), .C0(N430), .Y(N434) );
  OAI32X1TF U665 ( .A0(N202), .A1(REG_B[1]), .A2(N224), .B0(N592), .B1(N202), 
        .Y(N439) );
  OAI211X1TF U666 ( .A0(N1084), .A1(N120), .B0(N1063), .C0(N1062), .Y(N5060)
         );
  AOI22X1TF U667 ( .A0(IO_DATAINA[5]), .A1(N1159), .B0(N1170), .B1(N1074), .Y(
        N1062) );
  AOI22X1TF U668 ( .A0(IO_DATAINB[5]), .A1(N135), .B0(D_ADDR[6]), .B1(N1144), 
        .Y(N1063) );
  OAI211X1TF U669 ( .A0(N1084), .A1(N1143), .B0(N1083), .C0(N1082), .Y(N5150)
         );
  AOI22X1TF U670 ( .A0(IO_DATAINA[4]), .A1(N169), .B0(N1172), .B1(N1081), .Y(
        N1082) );
  AOI221X1TF U671 ( .A0(N221), .A1(N249), .B0(REG_A[3]), .B1(N166), .C0(N593), 
        .Y(N594) );
  OAI31X1TF U672 ( .A0(N748), .A1(N181), .A2(N801), .B0(N788), .Y(N593) );
  OAI21X1TF U673 ( .A0(REG_B[3]), .A1(N224), .B0(N592), .Y(N595) );
  AOI22X1TF U674 ( .A0(N796), .A1(N793), .B0(N703), .B1(N795), .Y(N597) );
  OAI211X1TF U675 ( .A0(N212), .A1(N119), .B0(N5850), .C0(N5840), .Y(N586) );
  AOI22X1TF U676 ( .A0(IO_DATAINB[4]), .A1(N135), .B0(D_ADDR[5]), .B1(N1144), 
        .Y(N1083) );
  INVX2TF U677 ( .A(N1061), .Y(N1084) );
  OAI211X1TF U678 ( .A0(N183), .A1(N710), .B0(N709), .C0(N708), .Y(N1061) );
  OAI21X1TF U679 ( .A0(N705), .A1(N775), .B0(N704), .Y(N706) );
  AOI22X1TF U680 ( .A0(N796), .A1(N737), .B0(N703), .B1(N766), .Y(N704) );
  INVX2TF U681 ( .A(N800), .Y(N703) );
  OAI22X1TF U682 ( .A0(N621), .A1(N209), .B0(N735), .B1(N773), .Y(N707) );
  OAI211X1TF U683 ( .A0(N1077), .A1(N120), .B0(N1057), .C0(N1056), .Y(N5030)
         );
  AOI22X1TF U684 ( .A0(IO_DATAINA[7]), .A1(N169), .B0(N1170), .B1(N1067), .Y(
        N1056) );
  OAI211X1TF U685 ( .A0(N186), .A1(N808), .B0(N807), .C0(N806), .Y(N1067) );
  OAI21X1TF U686 ( .A0(N801), .A1(N800), .B0(N799), .Y(N802) );
  AOI22X1TF U687 ( .A0(N798), .A1(N797), .B0(N796), .B1(N795), .Y(N799) );
  INVX2TF U688 ( .A(N591), .Y(N795) );
  OAI22X1TF U689 ( .A0(N245), .A1(N204), .B0(N752), .B1(N211), .Y(N520) );
  AOI22X1TF U690 ( .A0(IO_DATAINB[7]), .A1(N135), .B0(D_ADDR[8]), .B1(N1144), 
        .Y(N1057) );
  OAI211X1TF U691 ( .A0(N1077), .A1(N1143), .B0(N1076), .C0(N1075), .Y(N5120)
         );
  AOI22X1TF U692 ( .A0(IO_DATAINA[6]), .A1(N169), .B0(N1172), .B1(N1074), .Y(
        N1075) );
  OAI211X1TF U693 ( .A0(N184), .A1(N734), .B0(N733), .C0(N732), .Y(N1074) );
  AOI211X1TF U694 ( .A0(N796), .A1(N731), .B0(N730), .C0(N729), .Y(N732) );
  OAI22X1TF U695 ( .A0(N758), .A1(N800), .B0(N757), .B1(N728), .Y(N729) );
  AOI22X1TF U696 ( .A0(IO_DATAINB[6]), .A1(N136), .B0(D_ADDR[7]), .B1(N139), 
        .Y(N1076) );
  INVX2TF U697 ( .A(N1055), .Y(N1077) );
  OAI211X1TF U698 ( .A0(N185), .A1(N722), .B0(N721), .C0(N720), .Y(N1055) );
  OAI31X1TF U699 ( .A0(N182), .A1(N748), .A2(N716), .B0(N715), .Y(N717) );
  AOI22X1TF U700 ( .A0(N798), .A1(N714), .B0(N796), .B1(N713), .Y(N715) );
  INVX2TF U701 ( .A(N532), .Y(N796) );
  OAI22X1TF U702 ( .A0(N193), .A1(N408), .B0(N407), .B1(N782), .Y(N409) );
  INVX2TF U703 ( .A(N441), .Y(N714) );
  AOI31X1TF U704 ( .A0(N573), .A1(N403), .A2(N568), .B0(N805), .Y(N411) );
  AOI32X1TF U705 ( .A0(N249), .A1(REG_A[14]), .A2(N193), .B0(N765), .B1(
        REG_A[14]), .Y(N413) );
  AOI32X1TF U706 ( .A0(N249), .A1(REG_A[0]), .A2(N1150), .B0(N745), .B1(
        REG_A[0]), .Y(N746) );
  AOI211X1TF U707 ( .A0(REG_B[0]), .A1(N744), .B0(N743), .C0(N742), .Y(N747)
         );
  AOI31X1TF U708 ( .A0(N741), .A1(N740), .A2(N739), .B0(N773), .Y(N743) );
  INVX2TF U709 ( .A(N735), .Y(N736) );
  NOR4X1TF U710 ( .A(N604), .B(N603), .C(N602), .D(N601), .Y(N735) );
  NOR2X1TF U711 ( .A(N600), .B(N209), .Y(N602) );
  INVX2TF U712 ( .A(N622), .Y(N737) );
  NOR4BX1TF U713 ( .AN(N568), .B(N567), .C(N566), .D(N768), .Y(N622) );
  OAI32X4TF U714 ( .A0(N139), .A1(CODE_TYPE[4]), .A2(N203), .B0(N895), .B1(
        N139), .Y(N1170) );
  INVX2TF U715 ( .A(N1166), .Y(N1163) );
  NOR2X1TF U716 ( .A(N752), .B(N211), .Y(N359) );
  NOR2X1TF U717 ( .A(N245), .B(N216), .Y(N422) );
  NOR2X1TF U718 ( .A(N24), .B(N204), .Y(N360) );
  AOI32X1TF U719 ( .A0(N249), .A1(REG_A[15]), .A2(N194), .B0(N745), .B1(
        REG_A[15]), .Y(N362) );
  OAI21X1TF U720 ( .A0(N805), .A1(N600), .B0(N592), .Y(N745) );
  OAI211X1TF U721 ( .A0(N206), .A1(N245), .B0(N353), .C0(N430), .Y(N797) );
  OAI211X1TF U722 ( .A0(N189), .A1(N400), .B0(N399), .C0(N398), .Y(N401) );
  NOR2X1TF U723 ( .A(N24), .B(N213), .Y(N567) );
  NOR2X1TF U724 ( .A(N245), .B(N218), .Y(N604) );
  OAI22X1TF U725 ( .A0(N441), .A1(N576), .B0(N489), .B1(N396), .Y(N402) );
  AOI22X1TF U726 ( .A0(REG_B[2]), .A1(N404), .B0(N713), .B1(N181), .Y(N489) );
  OAI211X1TF U727 ( .A0(N245), .A1(N211), .B0(N395), .C0(N767), .Y(N713) );
  AOI221X1TF U728 ( .A0(REG_B[0]), .A1(N210), .B0(N1150), .B1(N204), .C0(
        REG_B[1]), .Y(N404) );
  OAI22X1TF U729 ( .A0(N24), .A1(N202), .B0(N752), .B1(N206), .Y(N394) );
  NOR2X1TF U730 ( .A(N24), .B(N217), .Y(N603) );
  OAI21X1TF U731 ( .A0(N1162), .A1(N1161), .B0(N1160), .Y(N1168) );
  OAI22X1TF U732 ( .A0(N191), .A1(N784), .B0(N783), .B1(N782), .Y(N785) );
  NOR2X1TF U733 ( .A(N752), .B(N212), .Y(N601) );
  NOR2X1TF U734 ( .A(N600), .B(N215), .Y(N566) );
  INVX2TF U735 ( .A(N775), .Y(N778) );
  NOR2X1TF U736 ( .A(N181), .B(N182), .Y(N779) );
  NOR2X2TF U737 ( .A(REG_B[2]), .B(N182), .Y(N780) );
  OAI211X1TF U738 ( .A0(N202), .A1(N245), .B0(N571), .C0(N570), .Y(N781) );
  OAI211X1TF U739 ( .A0(N774), .A1(N773), .B0(N772), .C0(N771), .Y(N786) );
  NOR2X1TF U740 ( .A(N214), .B(N752), .Y(N768) );
  NOR2X1TF U741 ( .A(N245), .B(N213), .Y(N770) );
  INVX2TF U742 ( .A(N766), .Y(N774) );
  OAI211X1TF U743 ( .A0(N210), .A1(N245), .B0(N574), .C0(N573), .Y(N766) );
  INVX2TF U744 ( .A(N224), .Y(N250) );
  OAI211X1TF U745 ( .A0(N192), .A1(N762), .B0(N761), .C0(N760), .Y(N763) );
  AOI32X1TF U746 ( .A0(N249), .A1(REG_A[13]), .A2(N192), .B0(N765), .B1(
        REG_A[13]), .Y(N760) );
  INVX2TF U747 ( .A(N224), .Y(N249) );
  OAI22X1TF U748 ( .A0(N758), .A1(N773), .B0(N757), .B1(N756), .Y(N759) );
  AOI22X1TF U749 ( .A0(REG_B[2]), .A1(N727), .B0(N726), .B1(N181), .Y(N757) );
  OAI211X1TF U750 ( .A0(N219), .A1(N245), .B0(N553), .C0(N5840), .Y(N726) );
  AOI221X1TF U751 ( .A0(N1150), .A1(N202), .B0(REG_B[0]), .B1(N206), .C0(
        REG_B[1]), .Y(N727) );
  INVX2TF U752 ( .A(N792), .Y(N773) );
  INVX2TF U753 ( .A(N725), .Y(N758) );
  OAI21X1TF U754 ( .A0(N752), .A1(N210), .B0(N428), .Y(N725) );
  INVX2TF U755 ( .A(N256), .Y(N350) );
  NOR2X1TF U756 ( .A(N860), .B(N854), .Y(N256) );
  NOR2X1TF U757 ( .A(N205), .B(N349), .Y(N852) );
  OR2X2TF U758 ( .A(N857), .B(N354), .Y(N868) );
  INVX2TF U759 ( .A(N855), .Y(N354) );
  INVX2TF U760 ( .A(N893), .Y(N358) );
  INVX2TF U761 ( .A(N224), .Y(N248) );
  OR2X2TF U762 ( .A(N860), .B(N261), .Y(N224) );
  INVX2TF U763 ( .A(N366), .Y(N261) );
  INVX2TF U764 ( .A(N705), .Y(N798) );
  NOR2X2TF U765 ( .A(N181), .B(REG_B[3]), .Y(N776) );
  INVX2TF U766 ( .A(N782), .Y(N755) );
  NOR2X4TF U767 ( .A(REG_B[0]), .B(REG_B[1]), .Y(N572) );
  AOI211X1TF U768 ( .A0(REG_A[11]), .A1(N153), .B0(N751), .C0(N750), .Y(N754)
         );
  NOR2X1TF U769 ( .A(N214), .B(N245), .Y(N750) );
  NOR2X2TF U770 ( .A(N1150), .B(N1124), .Y(N548) );
  NOR2X1TF U771 ( .A(N24), .B(N216), .Y(N751) );
  INVX2TF U772 ( .A(REG_B[1]), .Y(N1124) );
  OAI22X1TF U773 ( .A0(N254), .A1(N860), .B0(N892), .B1(N347), .Y(N790) );
  NAND2X2TF U774 ( .A(CODE_TYPE[3]), .B(N205), .Y(N860) );
  AOI21X1TF U775 ( .A0(N893), .A1(N26), .B0(N858), .Y(N254) );
  AOI22X1TF U776 ( .A0(N169), .A1(IO_DATAINA[0]), .B0(IO_STATUS[0]), .B1(N1158), .Y(N1174) );
  NOR2X1TF U777 ( .A(N26), .B(N1129), .Y(N1158) );
  AOI22X1TF U778 ( .A0(IO_DATAINB[0]), .A1(N136), .B0(D_ADDR[1]), .B1(N1144), 
        .Y(N1175) );
  INVX2TF U779 ( .A(N894), .Y(N892) );
  OAI22X1TF U780 ( .A0(N140), .A1(N635), .B0(N170), .B1(N699), .Y(N877) );
  OAI22X1TF U781 ( .A0(N667), .A1(N146), .B0(N221), .B1(N144), .Y(N878) );
  OAI22X1TF U782 ( .A0(N140), .A1(N629), .B0(N1136), .B1(N693), .Y(N1085) );
  OAI22X1TF U783 ( .A0(N661), .A1(N145), .B0(N213), .B1(N143), .Y(N1086) );
  OAI22X1TF U784 ( .A0(N141), .A1(N630), .B0(N1136), .B1(N694), .Y(N1064) );
  OAI22X1TF U785 ( .A0(N662), .A1(N145), .B0(N215), .B1(N143), .Y(N1065) );
  OAI22X1TF U786 ( .A0(N141), .A1(N627), .B0(N1136), .B1(N691), .Y(N1115) );
  OAI22X1TF U787 ( .A0(N659), .A1(N145), .B0(N220), .B1(N143), .Y(N1116) );
  OAI22X1TF U788 ( .A0(N140), .A1(N628), .B0(N1136), .B1(N692), .Y(N1104) );
  OAI22X1TF U789 ( .A0(N660), .A1(N145), .B0(N214), .B1(N143), .Y(N1105) );
  OAI22X1TF U790 ( .A0(N141), .A1(N625), .B0(N1136), .B1(N689), .Y(N1110) );
  OAI22X1TF U791 ( .A0(N657), .A1(N145), .B0(N211), .B1(N143), .Y(N1111) );
  OAI22X1TF U792 ( .A0(N140), .A1(N637), .B0(N1136), .B1(N701), .Y(N910) );
  OAI22X1TF U793 ( .A0(N669), .A1(N145), .B0(N202), .B1(N144), .Y(N911) );
  OAI22X1TF U794 ( .A0(N141), .A1(N633), .B0(N1136), .B1(N697), .Y(N1058) );
  OAI22X1TF U795 ( .A0(N665), .A1(N145), .B0(N217), .B1(N144), .Y(N1059) );
  OAI22X1TF U796 ( .A0(N141), .A1(N624), .B0(N1136), .B1(N688), .Y(N1121) );
  OAI22X1TF U797 ( .A0(N656), .A1(N146), .B0(N204), .B1(N144), .Y(N1122) );
  OAI22X1TF U798 ( .A0(N140), .A1(N634), .B0(N170), .B1(N698), .Y(N1078) );
  OAI22X1TF U799 ( .A0(N666), .A1(N146), .B0(N209), .B1(N143), .Y(N1079) );
  OAI22X1TF U800 ( .A0(N141), .A1(N631), .B0(N170), .B1(N695), .Y(N900) );
  OAI22X1TF U801 ( .A0(N663), .A1(N146), .B0(N218), .B1(N144), .Y(N901) );
  OAI22X1TF U802 ( .A0(N140), .A1(N632), .B0(N170), .B1(N696), .Y(N1071) );
  OAI22X1TF U803 ( .A0(N664), .A1(N146), .B0(N212), .B1(N143), .Y(N1072) );
  OAI22X1TF U804 ( .A0(N141), .A1(N623), .B0(N170), .B1(N687), .Y(N1138) );
  OAI22X1TF U805 ( .A0(N655), .A1(N146), .B0(N210), .B1(N144), .Y(N1139) );
  OAI22X1TF U806 ( .A0(N140), .A1(N626), .B0(N170), .B1(N690), .Y(N1099) );
  OAI22X1TF U807 ( .A0(N658), .A1(N146), .B0(N216), .B1(N144), .Y(N1100) );
  OAI22X1TF U808 ( .A0(N140), .A1(N636), .B0(N170), .B1(N700), .Y(N913) );
  OAI22X1TF U809 ( .A0(N668), .A1(N146), .B0(N219), .B1(N144), .Y(N914) );
  OAI22X1TF U810 ( .A0(N141), .A1(N638), .B0(N1136), .B1(N702), .Y(N907) );
  OAI22X1TF U811 ( .A0(N670), .A1(N145), .B0(N206), .B1(N143), .Y(N908) );
  AOI211X1TF U812 ( .A0(N468), .A1(N149), .B0(N517), .C0(N5140), .Y(N1096) );
  AOI211X1TF U813 ( .A0(N133), .A1(N753), .B0(N557), .C0(N556), .Y(N559) );
  AOI21X1TF U814 ( .A0(N250), .A1(N188), .B0(N127), .Y(N552) );
  AOI22X1TF U815 ( .A0(N509), .A1(N171), .B0(N475), .B1(N149), .Y(N560) );
  AOI221X1TF U816 ( .A0(N248), .A1(N213), .B0(N166), .B1(REG_A[9]), .C0(N138), 
        .Y(N561) );
  AOI211X1TF U817 ( .A0(N133), .A1(N541), .B0(N538), .C0(N535), .Y(N544) );
  AOI21X1TF U818 ( .A0(N250), .A1(N190), .B0(N127), .Y(N523) );
  AOI22X1TF U819 ( .A0(N511), .A1(N171), .B0(N477), .B1(N149), .Y(N546) );
  AOI221X1TF U820 ( .A0(N248), .A1(N220), .B0(N166), .B1(REG_A[11]), .C0(N138), 
        .Y(N547) );
  AOI211X1TF U821 ( .A0(N133), .A1(N777), .B0(N578), .C0(N577), .Y(N580) );
  AOI21X1TF U822 ( .A0(N250), .A1(N187), .B0(N127), .Y(N569) );
  AOI22X1TF U823 ( .A0(N508), .A1(N171), .B0(N474), .B1(N149), .Y(N581) );
  AOI221X1TF U824 ( .A0(N248), .A1(N215), .B0(N166), .B1(REG_A[8]), .C0(N138), 
        .Y(N583) );
  AOI22X1TF U825 ( .A0(N501), .A1(N244), .B0(N467), .B1(N148), .Y(N436) );
  AOI22X1TF U826 ( .A0(N133), .A1(N797), .B0(N792), .B1(N586), .Y(N598) );
  AOI22X1TF U827 ( .A0(N503), .A1(N244), .B0(N469), .B1(N148), .Y(N599) );
  AOI211X1TF U828 ( .A0(N133), .A1(N781), .B0(N707), .C0(N706), .Y(N708) );
  AOI21X1TF U829 ( .A0(N249), .A1(N183), .B0(N127), .Y(N621) );
  AOI22X1TF U830 ( .A0(N504), .A1(N171), .B0(N470), .B1(N149), .Y(N709) );
  AOI221X1TF U831 ( .A0(N249), .A1(N209), .B0(N166), .B1(REG_A[4]), .C0(N138), 
        .Y(N710) );
  AOI211X1TF U832 ( .A0(N133), .A1(N804), .B0(N803), .C0(N802), .Y(N806) );
  AOI211X1TF U833 ( .A0(REG_A[11]), .A1(N173), .B0(N751), .C0(N520), .Y(N591)
         );
  AOI21X1TF U834 ( .A0(N249), .A1(N186), .B0(N127), .Y(N794) );
  AOI22X1TF U835 ( .A0(N507), .A1(N244), .B0(N473), .B1(N149), .Y(N807) );
  AOI221X1TF U836 ( .A0(N248), .A1(N218), .B0(N166), .B1(REG_A[7]), .C0(N138), 
        .Y(N808) );
  AOI21X1TF U837 ( .A0(N250), .A1(N184), .B0(N127), .Y(N724) );
  AOI22X1TF U838 ( .A0(N505), .A1(N171), .B0(N471), .B1(N149), .Y(N733) );
  AOI221X1TF U839 ( .A0(N248), .A1(N217), .B0(N166), .B1(REG_A[5]), .C0(N138), 
        .Y(N734) );
  AOI211X1TF U840 ( .A0(N133), .A1(N719), .B0(N718), .C0(N717), .Y(N720) );
  AOI21X1TF U841 ( .A0(N250), .A1(N185), .B0(N127), .Y(N712) );
  AOI22X1TF U842 ( .A0(N506), .A1(N171), .B0(N472), .B1(N149), .Y(N721) );
  AOI221X1TF U843 ( .A0(N248), .A1(N212), .B0(N166), .B1(REG_A[6]), .C0(N138), 
        .Y(N722) );
  AOI221X1TF U844 ( .A0(N248), .A1(N204), .B0(N166), .B1(REG_A[14]), .C0(N138), 
        .Y(N408) );
  OAI31X1TF U845 ( .A0(N360), .A1(N422), .A2(N359), .B0(N133), .Y(N361) );
  AOI21X1TF U846 ( .A0(N572), .A1(N792), .B0(N126), .Y(N592) );
  AOI221X1TF U847 ( .A0(N248), .A1(N210), .B0(N166), .B1(REG_A[15]), .C0(N137), 
        .Y(N356) );
  AOI22X1TF U848 ( .A0(N572), .A1(REG_A[3]), .B0(N153), .B1(REG_A[1]), .Y(N353) );
  AOI22X1TF U849 ( .A0(N510), .A1(N244), .B0(N476), .B1(N148), .Y(N398) );
  AOI22X1TF U850 ( .A0(REG_A[10]), .A1(N397), .B0(N132), .B1(N406), .Y(N399)
         );
  AOI221X1TF U851 ( .A0(N789), .A1(REG_A[10]), .B0(N249), .B1(N214), .C0(N137), 
        .Y(N400) );
  AOI22X1TF U852 ( .A0(REG_A[10]), .A1(N173), .B0(N153), .B1(REG_A[12]), .Y(
        N395) );
  INVX2TF U853 ( .A(N572), .Y(N600) );
  AOI22X1TF U854 ( .A0(N572), .A1(REG_A[4]), .B0(N152), .B1(REG_A[2]), .Y(N571) );
  AOI221X1TF U855 ( .A0(N248), .A1(N216), .B0(N789), .B1(REG_A[12]), .C0(N137), 
        .Y(N784) );
  OAI31X1TF U856 ( .A0(N770), .A1(N769), .A2(N768), .B0(N132), .Y(N771) );
  AOI22X1TF U857 ( .A0(N512), .A1(N244), .B0(N478), .B1(N148), .Y(N772) );
  AOI22X1TF U858 ( .A0(N173), .A1(REG_A[12]), .B0(N153), .B1(REG_A[14]), .Y(
        N574) );
  AOI22X1TF U859 ( .A0(N572), .A1(REG_A[5]), .B0(N152), .B1(REG_A[3]), .Y(N553) );
  AOI221X1TF U860 ( .A0(N248), .A1(N211), .B0(N789), .B1(REG_A[13]), .C0(N137), 
        .Y(N762) );
  INVX2TF U861 ( .A(N1141), .Y(N1172) );
  NAND2X1TF U862 ( .A(OPER3_R3[1]), .B(N373), .Y(N1151) );
  NAND2X1TF U863 ( .A(OPER3_R3[0]), .B(N370), .Y(N1147) );
  OAI221XLTF U864 ( .A0(N579), .A1(NF), .B0(N203), .B1(N234), .C0(CODE_TYPE[2]), .Y(N258) );
  OAI2BB2XLTF U865 ( .B0(N754), .B1(N805), .A0N(N753), .A1N(N798), .Y(N764) );
  NAND2X1TF U866 ( .A(N755), .B(N776), .Y(N705) );
  CLKBUFX2TF U867 ( .A(N1151), .Y(N247) );
  CLKBUFX2TF U868 ( .A(N1147), .Y(N246) );
  INVX2TF U869 ( .A(N859), .Y(N881) );
  NAND2X1TF U870 ( .A(N562), .B(N1049), .Y(N335) );
  NOR4XLTF U871 ( .A(N27), .B(N882), .C(N881), .D(N273), .Y(N163) );
  NAND3X1TF U872 ( .A(I_ADDR[1]), .B(I_ADDR[2]), .C(I_ADDR[3]), .Y(N318) );
  NAND2X1TF U873 ( .A(N321), .B(I_ADDR[5]), .Y(N324) );
  NOR2BX1TF U874 ( .AN(N334), .B(N333), .Y(N164) );
  NAND2X1TF U875 ( .A(N861), .B(N208), .Y(N347) );
  NAND2X1TF U876 ( .A(N134), .B(N225), .Y(N854) );
  NOR4XLTF U877 ( .A(N564), .B(STATE[1]), .C(N226), .D(N257), .Y(N612) );
  NAND3X1TF U878 ( .A(N906), .B(N346), .C(START), .Y(N264) );
  NAND2X1TF U879 ( .A(N128), .B(N265), .Y(N323) );
  AOI2BB2X1TF U880 ( .B0(I_ADDR[1]), .B1(N322), .A0N(N328), .A1N(I_ADDR[1]), 
        .Y(N266) );
  NAND2X1TF U881 ( .A(N327), .B(N233), .Y(N267) );
  NAND4X1TF U882 ( .A(N1144), .B(N274), .C(N340), .D(N269), .Y(N1016) );
  NAND2X1TF U883 ( .A(I_ADDR[1]), .B(I_ADDR[2]), .Y(N317) );
  NAND4X1TF U884 ( .A(N682), .B(N681), .C(N680), .D(N679), .Y(N337) );
  NAND2BX1TF U885 ( .AN(N854), .B(N579), .Y(N857) );
  NAND2X1TF U886 ( .A(N159), .B(REG_A[6]), .Y(N425) );
  NAND2X1TF U887 ( .A(REG_A[7]), .B(N173), .Y(N589) );
  NAND4X1TF U888 ( .A(N425), .B(N351), .C(N5850), .D(N589), .Y(N804) );
  NAND2X1TF U889 ( .A(REG_A[10]), .B(N159), .Y(N419) );
  NAND2X1TF U890 ( .A(N548), .B(REG_A[8]), .Y(N426) );
  NAND2X1TF U891 ( .A(REG_A[9]), .B(N153), .Y(N588) );
  NAND4X1TF U892 ( .A(N419), .B(N426), .C(N352), .D(N588), .Y(N541) );
  NAND2X1TF U893 ( .A(N159), .B(REG_A[2]), .Y(N430) );
  AOI222XLTF U894 ( .A0(N804), .A1(N780), .B0(N541), .B1(N776), .C0(N797), 
        .C1(N779), .Y(N357) );
  OA22X1TF U895 ( .A0(N357), .A1(N782), .B0(N194), .B1(N356), .Y(N363) );
  AO21X1TF U896 ( .A0(N820), .A1(N367), .B0(N880), .Y(N1145) );
  NAND2X1TF U897 ( .A(N548), .B(REG_A[3]), .Y(N740) );
  NAND2X1TF U898 ( .A(N755), .B(N780), .Y(N576) );
  NAND2X1TF U899 ( .A(N159), .B(REG_A[11]), .Y(N767) );
  AO21X1TF U900 ( .A0(N189), .A1(N250), .B0(N127), .Y(N397) );
  AO21X1TF U901 ( .A0(N132), .A1(N173), .B0(N126), .Y(N765) );
  NAND2X1TF U902 ( .A(N159), .B(REG_A[13]), .Y(N573) );
  NAND2X1TF U903 ( .A(N153), .B(REG_A[12]), .Y(N403) );
  NAND2X1TF U904 ( .A(N548), .B(REG_A[11]), .Y(N568) );
  NAND2X1TF U905 ( .A(N404), .B(N181), .Y(N716) );
  AOI222XLTF U906 ( .A0(N719), .A1(N780), .B0(N406), .B1(N776), .C0(N714), 
        .C1(N779), .Y(N407) );
  OAI221XLTF U907 ( .A0(REG_A[1]), .A1(N224), .B0(N202), .B1(N738), .C0(N788), 
        .Y(N440) );
  NAND2X1TF U908 ( .A(REG_A[9]), .B(N572), .Y(N551) );
  NAND2X1TF U909 ( .A(REG_A[7]), .B(N152), .Y(N550) );
  NAND4X1TF U910 ( .A(N427), .B(N550), .C(N426), .D(N425), .Y(N723) );
  AOI222XLTF U911 ( .A0(N731), .A1(N780), .B0(N723), .B1(N776), .C0(N725), 
        .C1(N779), .Y(N437) );
  NAND2X1TF U912 ( .A(N182), .B(N755), .Y(N728) );
  NAND2X1TF U913 ( .A(N181), .B(N727), .Y(N555) );
  AOI2BB2X1TF U914 ( .B0(N792), .B1(N434), .A0N(N728), .A1N(N555), .Y(N435) );
  NAND2X1TF U915 ( .A(N158), .B(REG_A[3]), .Y(N570) );
  NAND2X1TF U916 ( .A(N548), .B(REG_A[5]), .Y(N565) );
  NAND2X1TF U917 ( .A(N590), .B(N776), .Y(N532) );
  NAND2X1TF U918 ( .A(REG_A[7]), .B(N158), .Y(N563) );
  NAND4BX1TF U919 ( .AN(N770), .B(N5000), .C(N491), .D(N563), .Y(N711) );
  OAI221XLTF U920 ( .A0(REG_A[2]), .A1(N224), .B0(N219), .B1(N738), .C0(N788), 
        .Y(N5020) );
  NAND2X1TF U921 ( .A(N159), .B(REG_A[8]), .Y(N587) );
  NAND4X1TF U922 ( .A(N551), .B(N550), .C(N549), .D(N587), .Y(N753) );
  OAI2BB2XLTF U923 ( .B0(N552), .B1(N213), .A0N(N731), .A1N(N792), .Y(N557) );
  NAND2X1TF U924 ( .A(N158), .B(REG_A[4]), .Y(N5840) );
  NAND4BBX1TF U925 ( .AN(N566), .BN(N601), .C(N565), .D(N563), .Y(N777) );
  NAND4BX1TF U926 ( .AN(N750), .B(N589), .C(N588), .D(N587), .Y(N793) );
  NAND2X1TF U927 ( .A(N590), .B(N780), .Y(N800) );
  AOI2BB2X1TF U928 ( .B0(REG_A[3]), .B1(N595), .A0N(N182), .A1N(N594), .Y(N596) );
  NAND4X1TF U929 ( .A(N599), .B(N598), .C(N597), .D(N596), .Y(N1081) );
  OAI2BB2XLTF U930 ( .B0(N712), .B1(N212), .A0N(N711), .A1N(N792), .Y(N718) );
  OAI2BB2XLTF U931 ( .B0(N724), .B1(N217), .A0N(N723), .A1N(N792), .Y(N730) );
  OAI221XLTF U932 ( .A0(REG_A[0]), .A1(N224), .B0(N206), .B1(N738), .C0(N788), 
        .Y(N744) );
  NAND2X1TF U933 ( .A(N159), .B(REG_A[1]), .Y(N741) );
  AO22X1TF U934 ( .A0(N500), .A1(N244), .B0(N466), .B1(N148), .Y(N742) );
  NAND2X1TF U935 ( .A(REG_B[3]), .B(N755), .Y(N756) );
  AO21X1TF U936 ( .A0(N250), .A1(N191), .B0(N765), .Y(N787) );
  AOI222XLTF U937 ( .A0(N781), .A1(N780), .B0(N779), .B1(N778), .C0(N777), 
        .C1(N776), .Y(N783) );
  OAI2BB2XLTF U938 ( .B0(N794), .B1(N218), .A0N(N793), .A1N(N792), .Y(N803) );
  NAND2X1TF U939 ( .A(N842), .B(N238), .Y(N826) );
  NAND2X1TF U940 ( .A(N842), .B(N236), .Y(N830) );
  NAND2X1TF U941 ( .A(N842), .B(N237), .Y(N840) );
  OAI2BB2XLTF U942 ( .B0(N861), .B1(N860), .A0N(N859), .A1N(N858), .Y(N863) );
  NAND2X1TF U943 ( .A(N869), .B(N415), .Y(N866) );
  OAI22X1TF U944 ( .A0(N416), .A1(N866), .B0(N884), .B1(N872), .Y(N898) );
  NAND3X1TF U945 ( .A(N130), .B(N894), .C(N893), .Y(N1129) );
  AO22X1TF U946 ( .A0(N917), .A1(N236), .B0(N916), .B1(I_DATAIN[6]), .Y(N4670)
         );
  AO22X1TF U947 ( .A0(N917), .A1(N237), .B0(N916), .B1(I_DATAIN[5]), .Y(N4680)
         );
  AO22X1TF U948 ( .A0(N917), .A1(N238), .B0(N916), .B1(I_DATAIN[4]), .Y(N4690)
         );
  AO22X1TF U949 ( .A0(N917), .A1(OPER3_R3[2]), .B0(N916), .B1(I_DATAIN[2]), 
        .Y(N4710) );
  AO22X1TF U950 ( .A0(N917), .A1(OPER3_R3[1]), .B0(N916), .B1(I_DATAIN[1]), 
        .Y(N4720) );
  AO22X1TF U951 ( .A0(N917), .A1(OPER3_R3[0]), .B0(N916), .B1(I_DATAIN[0]), 
        .Y(N4730) );
  AO22X1TF U952 ( .A0(N919), .A1(CF_BUF), .B0(N918), .B1(CF), .Y(N4740) );
  AO22X1TF U953 ( .A0(N1054), .A1(CODE_TYPE[3]), .B0(N1053), .B1(I_DATAIN[6]), 
        .Y(N493) );
  AO22X1TF U954 ( .A0(N1054), .A1(CODE_TYPE[2]), .B0(N1053), .B1(I_DATAIN[5]), 
        .Y(N494) );
  AO22X1TF U955 ( .A0(N1054), .A1(N27), .B0(N1053), .B1(I_DATAIN[4]), .Y(N495)
         );
  AO22X1TF U956 ( .A0(N1054), .A1(\OPER1_R1[2] ), .B0(N1053), .B1(I_DATAIN[2]), 
        .Y(N497) );
  AOI2BB2X1TF U957 ( .B0(N25), .B1(N1054), .A0N(N1054), .A1N(I_DATAIN[1]), .Y(
        N498) );
  AO22X1TF U958 ( .A0(N1054), .A1(N222), .B0(N1053), .B1(I_DATAIN[0]), .Y(N499) );
  AOI2BB2X1TF U959 ( .B0(IO_DATAINB[8]), .B1(N136), .A0N(N131), .A1N(N429), 
        .Y(N1069) );
  AOI2BB2X1TF U960 ( .B0(IO_DATAINB[9]), .B1(N136), .A0N(N131), .A1N(N424), 
        .Y(N1091) );
  AOI2BB2X1TF U961 ( .B0(IO_DATAINA[2]), .B1(N1159), .A0N(N1096), .A1N(N1143), 
        .Y(N1097) );
  AOI2BB2X1TF U962 ( .B0(IO_DATAINB[12]), .B1(N136), .A0N(N131), .A1N(N423), 
        .Y(N1103) );
  AOI2BB2X1TF U963 ( .B0(IO_DATAINB[10]), .B1(N136), .A0N(N131), .A1N(N421), 
        .Y(N1108) );
  AOI2BB2X1TF U964 ( .B0(IO_DATAINB[11]), .B1(N136), .A0N(N131), .A1N(N418), 
        .Y(N1120) );
endmodule


module SCPU_SRAM_8BIT_ALU_SPI_TOP_VG ( CLK, RST_N, CTRL_MODE, CTRL_BGN, CPU_BGN, 
        LOAD_N, CTRL_SI, ADC_PI, CTRL_RDY, CTRL_SO, NXT, SCLK1, SCLK2, LAT, 
        SPI_SO );
  input [1:0] CTRL_MODE;
  input [15:0] ADC_PI;
  output [1:0] NXT;
  input CLK, RST_N, CTRL_BGN, CPU_BGN, LOAD_N, CTRL_SI;
  output CTRL_RDY, CTRL_SO, SCLK1, SCLK2, LAT, SPI_SO;
  wire   CEN_AFTER_MUX, WEN_AFTER_MUX, I_CLK, I_RST_N, I_CTRL_BGN, I_CPU_BGN,
         I_LOAD_N, I_CTRL_SI, I_CTRL_SO, I_SCLK1, I_SCLK2, I_SPI_SO,
         SCPU_CTRL_SPI_CEN, \SCPU_CTRL_SPI_IO_DATAOUTB[0] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[1] , \SCPU_CTRL_SPI_IO_DATAOUTB[2] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[3] , \SCPU_CTRL_SPI_IO_DATAOUTB[4] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[5] , \SCPU_CTRL_SPI_IO_DATAOUTB[6] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[7] , \SCPU_CTRL_SPI_IO_DATAOUTB[8] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[9] , \SCPU_CTRL_SPI_IO_DATAOUTB[10] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[11] , \SCPU_CTRL_SPI_IO_DATAOUTB[12] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[0] , \SCPU_CTRL_SPI_IO_DATAOUTA[1] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[2] , \SCPU_CTRL_SPI_IO_DATAOUTA[3] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[4] , \SCPU_CTRL_SPI_IO_DATAOUTA[5] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[6] , \SCPU_CTRL_SPI_IO_DATAOUTA[7] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[8] , \SCPU_CTRL_SPI_IO_DATAOUTA[9] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[10] , \SCPU_CTRL_SPI_IO_DATAOUTA[11] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[12] , \SCPU_CTRL_SPI_IO_CONTROL[0] ,
         \SCPU_CTRL_SPI_IO_CONTROL[1] , \SCPU_CTRL_SPI_IO_CONTROL[2] ,
         \SCPU_CTRL_SPI_IO_CONTROL[3] , \SCPU_CTRL_SPI_IO_CONTROL[4] ,
         \SCPU_CTRL_SPI_IO_CONTROL[5] , \SCPU_CTRL_SPI_IO_CONTROL[6] ,
         SCPU_CTRL_SPI_D_WE, SCPU_CTRL_SPI_IS_I_ADDR, SCPU_CTRL_SPI_CCT_N54,
         SCPU_CTRL_SPI_CCT_N53, SCPU_CTRL_SPI_CCT_N51, SCPU_CTRL_SPI_CCT_N50,
         SCPU_CTRL_SPI_CCT_N49, SCPU_CTRL_SPI_CCT_N24,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] , \SCPU_CTRL_SPI_CCT_REG_BITS[1] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[2] , \SCPU_CTRL_SPI_CCT_REG_BITS[3] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[4] , \SCPU_CTRL_SPI_CCT_REG_BITS[5] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[6] , \SCPU_CTRL_SPI_CCT_REG_BITS[7] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[8] , \SCPU_CTRL_SPI_CCT_REG_BITS[9] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[10] , \SCPU_CTRL_SPI_CCT_REG_BITS[11] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[12] , \SCPU_CTRL_SPI_CCT_REG_BITS[13] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[14] , \SCPU_CTRL_SPI_CCT_REG_BITS[15] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[16] , \SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ,
         SCPU_CTRL_SPI_PUT_N108, SCPU_CTRL_SPI_PUT_N107,
         SCPU_CTRL_SPI_PUT_N106, \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ,
         \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ,
         \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ,
         \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] , \SCPU_CTRL_SPI_PUT_SPI_STATE[0] ,
         \SCPU_CTRL_SPI_PUT_SPI_STATE[1] , \SCPU_CTRL_SPI_PUT_CNT_STATE[1] ,
         \SCPU_CTRL_SPI_PUT_CNT_STATE[2] , N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, N45, N78, N79, N80, N81, N82, N83,
         N84, N85, N86, N91, N93, N100, N102, N103, N158, N189, N190, N191,
         N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202,
         N203, N204, N205, N206, N207, N208, N209, N210, N212, N213, N214,
         N215, N216, N218, N219, N220, N221, N222, N233, N234, N241, N270,
         N271, N272, N273, N274, N275, N277, N278, N279, N280, N281, N282,
         N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293,
         N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304,
         N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315,
         N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326,
         N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337,
         N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, N348,
         N349, N350, N351, N352, N353, N354, N355, N356, N357, N358, N359,
         N360, N361, N362, N363, N364, N365, N366, N367, N368, N369, N370,
         N371, N372, N373, N374, N375, N376, N377, N378, N379, N380, N381,
         N382, N383, N384, N385, N386, N387, N388, N389, N390, N391, N392,
         N393, N394, N395, N396, N397, N398, N399, N400, N401, N402, N403,
         N404, N405, N406, N407, N408, N409, N410, N411, N412, N413, N414,
         N415, N416, N417, N418, N419, N420, N421, N422, N423, N424, N425,
         N426, N427, N428;
  wire   [8:0] A_AFTER_MUX;
  wire   [7:0] D_AFTER_MUX;
  wire   [7:0] Q_FROM_SRAM;
  wire   [1:0] I_CTRL_MODE;
  wire   [15:0] I_ADC_PI;
  wire   [1:0] I_NXT;
  wire   [8:0] SCPU_CTRL_SPI_A_SPI;
  wire   [12:0] SCPU_CTRL_SPI_POUT;
  wire   [12:0] SCPU_CTRL_SPI_FOUT;
  wire   [9:0] SCPU_CTRL_SPI_IO_OFFSET;
  wire   [15:0] SCPU_CTRL_SPI_IO_DATAINA;
  wire   [0:0] SCPU_CTRL_SPI_IO_STATUS;
  wire   [7:0] SCPU_CTRL_SPI_D_DATAOUT;
  wire   [8:1] SCPU_CTRL_SPI_D_ADDR;
  wire   [8:0] SCPU_CTRL_SPI_I_ADDR;
  wire   [7:0] SCPU_CTRL_SPI_D_DATAIN;
  wire   [7:0] SCPU_CTRL_SPI_I_DATAIN;
  wire   [7:1] SCPU_CTRL_SPI_PUT_SRAM_REGS;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21;

  RA1SHD_IBM512X8 sram ( .Q(Q_FROM_SRAM), .A(A_AFTER_MUX), .D(D_AFTER_MUX), 
        .CLK(I_CLK), .CEN(CEN_AFTER_MUX), .WEN(WEN_AFTER_MUX) );
  PIC ipad_clk ( .IE(1'b1), .P(CLK), .Y(I_CLK) );
  PIC ipad_rst_n ( .IE(1'b1), .P(RST_N), .Y(I_RST_N) );
  PIC ipad_ctrl_mode0 ( .IE(1'b1), .P(CTRL_MODE[0]), .Y(I_CTRL_MODE[0]) );
  PIC ipad_ctrl_mode1 ( .IE(1'b1), .P(CTRL_MODE[1]), .Y(I_CTRL_MODE[1]) );
  PIC ipad_ctrl_bgn ( .IE(1'b1), .P(CTRL_BGN), .Y(I_CTRL_BGN) );
  PIC ipad_cpu_str ( .IE(1'b1), .P(CPU_BGN), .Y(I_CPU_BGN) );
  PIC ipad_load_n ( .IE(1'b1), .P(LOAD_N), .Y(I_LOAD_N) );
  PIC ipad_ctrl_si ( .IE(1'b1), .P(CTRL_SI), .Y(I_CTRL_SI) );
  PIC ipad_adc_pi0 ( .IE(1'b1), .P(ADC_PI[0]), .Y(I_ADC_PI[0]) );
  PIC ipad_adc_pi1 ( .IE(1'b1), .P(ADC_PI[1]), .Y(I_ADC_PI[1]) );
  PIC ipad_adc_pi2 ( .IE(1'b1), .P(ADC_PI[2]), .Y(I_ADC_PI[2]) );
  PIC ipad_adc_pi3 ( .IE(1'b1), .P(ADC_PI[3]), .Y(I_ADC_PI[3]) );
  PIC ipad_adc_pi4 ( .IE(1'b1), .P(ADC_PI[4]), .Y(I_ADC_PI[4]) );
  PIC ipad_adc_pi5 ( .IE(1'b1), .P(ADC_PI[5]), .Y(I_ADC_PI[5]) );
  PIC ipad_adc_pi6 ( .IE(1'b1), .P(ADC_PI[6]), .Y(I_ADC_PI[6]) );
  PIC ipad_adc_pi7 ( .IE(1'b1), .P(ADC_PI[7]), .Y(I_ADC_PI[7]) );
  PIC ipad_adc_pi8 ( .IE(1'b1), .P(ADC_PI[8]), .Y(I_ADC_PI[8]) );
  PIC ipad_adc_pi9 ( .IE(1'b1), .P(ADC_PI[9]), .Y(I_ADC_PI[9]) );
  PIC ipad_adc_pi10 ( .IE(1'b1), .P(ADC_PI[10]), .Y(I_ADC_PI[10]) );
  PIC ipad_adc_pi11 ( .IE(1'b1), .P(ADC_PI[11]), .Y(I_ADC_PI[11]) );
  PIC ipad_adc_pi12 ( .IE(1'b1), .P(ADC_PI[12]), .Y(I_ADC_PI[12]) );
  PIC ipad_adc_pi13 ( .IE(1'b1), .P(ADC_PI[13]), .Y(I_ADC_PI[13]) );
  PIC ipad_adc_pi14 ( .IE(1'b1), .P(ADC_PI[14]), .Y(I_ADC_PI[14]) );
  PIC ipad_adc_pi15 ( .IE(1'b1), .P(ADC_PI[15]), .Y(I_ADC_PI[15]) );
  POC8B opad_ctrl_rdy ( .A(N220), .P(CTRL_RDY) );
  POC8B opad_ctrl_so ( .A(I_CTRL_SO), .P(CTRL_SO) );
  POC8B opad_nxt0 ( .A(I_NXT[0]), .P(NXT[0]) );
  POC8B opad_nxt1 ( .A(I_NXT[1]), .P(NXT[1]) );
  POC8B opad_sclk1 ( .A(I_SCLK1), .P(SCLK1) );
  POC8B opad_sclk2 ( .A(I_SCLK2), .P(SCLK2) );
  POC8B opad_lat ( .A(N222), .P(LAT) );
  POC8B opad_spi_so ( .A(I_SPI_SO), .P(SPI_SO) );
  SHARE_SUPERALU_VG \scpu_ctrl_spi/ALU_01  ( .CLK(I_CLK), .RST_N(I_RST_N), .X_IN(
        {\SCPU_CTRL_SPI_IO_DATAOUTA[12] , \SCPU_CTRL_SPI_IO_DATAOUTA[11] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[10] , \SCPU_CTRL_SPI_IO_DATAOUTA[9] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[8] , \SCPU_CTRL_SPI_IO_DATAOUTA[7] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[6] , \SCPU_CTRL_SPI_IO_DATAOUTA[5] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[4] , \SCPU_CTRL_SPI_IO_DATAOUTA[3] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[2] , \SCPU_CTRL_SPI_IO_DATAOUTA[1] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[0] }), .Y_IN({
        \SCPU_CTRL_SPI_IO_DATAOUTB[12] , \SCPU_CTRL_SPI_IO_DATAOUTB[11] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[10] , \SCPU_CTRL_SPI_IO_DATAOUTB[9] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[8] , \SCPU_CTRL_SPI_IO_DATAOUTB[7] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[6] , \SCPU_CTRL_SPI_IO_DATAOUTB[5] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[4] , \SCPU_CTRL_SPI_IO_DATAOUTB[3] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[2] , \SCPU_CTRL_SPI_IO_DATAOUTB[1] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[0] }), .ALU_START(N390), .ALU_TYPE({
        \SCPU_CTRL_SPI_IO_CONTROL[4] , \SCPU_CTRL_SPI_IO_CONTROL[3] , 
        \SCPU_CTRL_SPI_IO_CONTROL[2] }), .MODE_TYPE({
        \SCPU_CTRL_SPI_IO_CONTROL[1] , \SCPU_CTRL_SPI_IO_CONTROL[0] }), 
        .OFFSET(SCPU_CTRL_SPI_IO_OFFSET), .FOUT(SCPU_CTRL_SPI_FOUT), .POUT(
        SCPU_CTRL_SPI_POUT), .ALU_IS_DONE(SCPU_CTRL_SPI_IO_STATUS[0]) );
  SERIAL_CPU_8BIT_VG \scpu_ctrl_spi/uut  ( .CLK(I_CLK), .ENABLE(1'b0), .RST_N(
        I_RST_N), .START(I_CPU_BGN), .I_DATAIN(SCPU_CTRL_SPI_I_DATAIN), 
        .D_DATAIN(SCPU_CTRL_SPI_D_DATAIN), .IS_I_ADDR(SCPU_CTRL_SPI_IS_I_ADDR), 
        .NXT(I_NXT), .I_ADDR(SCPU_CTRL_SPI_I_ADDR), .D_ADDR({
        SCPU_CTRL_SPI_D_ADDR, SYNOPSYS_UNCONNECTED__0}), .D_WE(
        SCPU_CTRL_SPI_D_WE), .D_DATAOUT(SCPU_CTRL_SPI_D_DATAOUT), .IO_STATUS({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, N221, SCPU_CTRL_SPI_IO_STATUS[0]}), .IO_CONTROL({
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, \SCPU_CTRL_SPI_IO_CONTROL[6] , 
        \SCPU_CTRL_SPI_IO_CONTROL[5] , \SCPU_CTRL_SPI_IO_CONTROL[4] , 
        \SCPU_CTRL_SPI_IO_CONTROL[3] , \SCPU_CTRL_SPI_IO_CONTROL[2] , 
        \SCPU_CTRL_SPI_IO_CONTROL[1] , \SCPU_CTRL_SPI_IO_CONTROL[0] }), 
        .IO_DATAINA(SCPU_CTRL_SPI_IO_DATAINA), .IO_DATAINB({1'b0, 1'b0, 1'b0, 
        SCPU_CTRL_SPI_POUT}), .IO_DATAOUTA({SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        \SCPU_CTRL_SPI_IO_DATAOUTA[12] , \SCPU_CTRL_SPI_IO_DATAOUTA[11] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[10] , \SCPU_CTRL_SPI_IO_DATAOUTA[9] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[8] , \SCPU_CTRL_SPI_IO_DATAOUTA[7] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[6] , \SCPU_CTRL_SPI_IO_DATAOUTA[5] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[4] , \SCPU_CTRL_SPI_IO_DATAOUTA[3] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[2] , \SCPU_CTRL_SPI_IO_DATAOUTA[1] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[0] }), .IO_DATAOUTB({
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, \SCPU_CTRL_SPI_IO_DATAOUTB[12] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[11] , \SCPU_CTRL_SPI_IO_DATAOUTB[10] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[9] , \SCPU_CTRL_SPI_IO_DATAOUTB[8] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[7] , \SCPU_CTRL_SPI_IO_DATAOUTB[6] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[5] , \SCPU_CTRL_SPI_IO_DATAOUTB[4] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[3] , \SCPU_CTRL_SPI_IO_DATAOUTB[2] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[1] , \SCPU_CTRL_SPI_IO_DATAOUTB[0] }), 
        .IO_OFFSET({SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SCPU_CTRL_SPI_IO_OFFSET}) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[5]  ( .D(N158), .RN(
        SCPU_CTRL_SPI_CCT_N53), .CK(I_CLK), .QN(N286) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[3]  ( .D(N158), .RN(
        SCPU_CTRL_SPI_CCT_N51), .CK(I_CLK), .QN(N285) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[2]  ( .D(N158), .RN(
        SCPU_CTRL_SPI_CCT_N50), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[1]  ( .D(N158), .RN(
        SCPU_CTRL_SPI_CCT_N49), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[6]  ( .D(N158), .RN(
        SCPU_CTRL_SPI_CCT_N54), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[4]  ( .D(N45), .CK(I_CLK), 
        .SN(N44), .RN(N43), .QN(N282) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[0]  ( .D(N33), .CK(I_CLK), 
        .SN(N32), .RN(N31), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .QN(N281)
         );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[3]  ( .D(N42), .CK(I_CLK), 
        .SN(N41), .RN(N40), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] ), .QN(N279)
         );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[2]  ( .D(N39), .CK(I_CLK), 
        .SN(N38), .RN(N37), .QN(N278) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[1]  ( .D(N36), .CK(I_CLK), 
        .SN(N35), .RN(N34), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ), .QN(N277)
         );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[7]  ( .D(N204), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[7]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[6]  ( .D(N198), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[6]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[5]  ( .D(N199), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[5]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[4]  ( .D(N200), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[4]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[3]  ( .D(N201), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[3]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[2]  ( .D(N202), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[2]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[1]  ( .D(N203), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[1]) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[7]  ( .D(N189), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[7] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[6]  ( .D(N190), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[6] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[5]  ( .D(N191), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[5] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[4]  ( .D(N192), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[4] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[3]  ( .D(N193), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[3] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[2]  ( .D(N194), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[2] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[1]  ( .D(N195), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[1] ) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[0]  ( .D(N197), .CK(I_CLK), .Q(
        I_SPI_SO) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[0]  ( .D(N196), .CK(I_CLK), .Q(
        I_CTRL_SO) );
  DFFQX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[4]  ( .D(N215), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ) );
  DFFSX2TF \scpu_ctrl_spi/put/cnt_state_reg[0]  ( .D(SCPU_CTRL_SPI_PUT_N106), 
        .CK(I_CLK), .SN(N271), .Q(N288), .QN(N102) );
  DFFQX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[0]  ( .D(N214), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ) );
  DFFRX1TF \scpu_ctrl_spi/put/spi_state_reg[0]  ( .D(N209), .CK(I_CLK), .RN(
        N271), .Q(\SCPU_CTRL_SPI_PUT_SPI_STATE[0] ) );
  DFFRX1TF \scpu_ctrl_spi/put/cnt_state_reg[1]  ( .D(SCPU_CTRL_SPI_PUT_N107), 
        .CK(I_CLK), .RN(N271), .Q(\SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .QN(N284)
         );
  DFFNSRX4TF \scpu_ctrl_spi/put/spi_MUX_reg  ( .D(N213), .CKN(I_CLK), .SN(1'b1), .RN(1'b1), .Q(N301), .QN(N103) );
  DFFNSRXLTF \scpu_ctrl_spi/cct/D_WE_reg  ( .D(N218), .CKN(I_CLK), .SN(1'b1), 
        .RN(1'b1), .QN(N93) );
  DFFNSRX1TF \scpu_ctrl_spi/put/sram_addr_reg[7]  ( .D(N85), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[7]), .QN(N289) );
  DFFNSRXLTF \scpu_ctrl_spi/cct/CEN_reg  ( .D(N219), .CKN(I_CLK), .SN(1'b1), 
        .RN(1'b1), .Q(SCPU_CTRL_SPI_CEN) );
  DFFNSRXLTF \scpu_ctrl_spi/put/sram_addr_reg[8]  ( .D(N86), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[8]) );
  DFFQX1TF \scpu_ctrl_spi/cct/ctrl_state_reg[0]  ( .D(N216), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ) );
  EDFFTRXLTF \scpu_ctrl_spi/cct/ctrl_state_reg[1]  ( .RN(I_CTRL_BGN), .D(1'b1), 
        .E(N234), .CK(I_CLK), .Q(N283), .QN(N91) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[16]  ( .D(I_CTRL_SI), .E(N241), 
        .CK(I_CLK), .Q(\SCPU_CTRL_SPI_CCT_REG_BITS[16] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[15]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[16] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[15] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[14]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[15] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[14] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[13]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[14] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[13] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[12]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[13] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[12] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[11]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[12] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[11] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[10]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[11] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[10] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[9]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[10] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[9] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[8]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[9] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[8] ) );
  DFFRX2TF \scpu_ctrl_spi/put/spi_state_reg[2]  ( .D(N212), .CK(I_CLK), .RN(
        N270), .Q(N287), .QN(N100) );
  DFFRX2TF \scpu_ctrl_spi/put/spi_state_reg[1]  ( .D(N210), .CK(I_CLK), .RN(
        N270), .Q(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .QN(N280) );
  DFFRX2TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[0]  ( .D(N205), .CK(I_CLK), 
        .RN(N271), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .QN(N290) );
  DFFRX2TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[3]  ( .D(N208), .CK(I_CLK), 
        .RN(N271), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ), .QN(N292) );
  DFFRX1TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[1]  ( .D(N206), .CK(I_CLK), 
        .RN(N270), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ) );
  DFFRX1TF \scpu_ctrl_spi/put/cnt_state_reg[2]  ( .D(SCPU_CTRL_SPI_PUT_N108), 
        .CK(I_CLK), .RN(N270), .Q(\SCPU_CTRL_SPI_PUT_CNT_STATE[2] ) );
  DFFRX1TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[2]  ( .D(N207), .CK(I_CLK), 
        .RN(N270), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[1]  ( .D(N79), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[1]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[3]  ( .D(N81), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[3]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[5]  ( .D(N83), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[5]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[2]  ( .D(N80), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[2]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[6]  ( .D(N84), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[6]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[4]  ( .D(N82), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[4]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[0]  ( .D(N78), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[0]), .QN(N291) );
  OR2X2TF U246 ( .A(SCPU_CTRL_SPI_IS_I_ADDR), .B(I_CTRL_BGN), .Y(N380) );
  CLKBUFX2TF U247 ( .A(N422), .Y(N294) );
  CLKBUFX2TF U248 ( .A(N422), .Y(N295) );
  INVX2TF U249 ( .A(N270), .Y(N422) );
  CLKBUFX2TF U250 ( .A(\SCPU_CTRL_SPI_IO_CONTROL[6] ), .Y(N270) );
  NOR3X1TF U251 ( .A(\SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .B(N102), .C(N103), 
        .Y(I_SCLK2) );
  NOR2BX1TF U252 ( .AN(I_ADC_PI[15]), .B(N390), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[15]) );
  NOR2BX1TF U253 ( .AN(I_ADC_PI[14]), .B(N390), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[14]) );
  AO21X1TF U254 ( .A0(N277), .A1(N424), .B0(N278), .Y(N233) );
  OAI21X1TF U255 ( .A0(N426), .A1(N427), .B0(N233), .Y(N39) );
  INVX2TF U256 ( .A(N299), .Y(N368) );
  OA21XLTF U257 ( .A0(\SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .A1(I_CTRL_MODE[0]), 
        .B0(N323), .Y(N234) );
  CLKBUFX2TF U258 ( .A(SCPU_CTRL_SPI_CCT_N24), .Y(N241) );
  AO21XLTF U272 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ), .A1(N296), .B0(
        N297), .Y(SCPU_CTRL_SPI_CCT_N50) );
  OR2X1TF U273 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ), .B(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .Y(N296) );
  OAI21XLTF U274 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .A1(N330), .B0(
        N329), .Y(N214) );
  NOR3X1TF U275 ( .A(N299), .B(N283), .C(N367), .Y(SCPU_CTRL_SPI_CCT_N24) );
  AO21XLTF U276 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ), .A1(N298), .B0(
        N299), .Y(SCPU_CTRL_SPI_CCT_N54) );
  AOI32X1TF U277 ( .A0(SCPU_CTRL_SPI_A_SPI[0]), .A1(N270), .A2(N426), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[0] ), .B1(N294), .Y(N420) );
  OAI21XLTF U278 ( .A0(N325), .A1(N286), .B0(N298), .Y(SCPU_CTRL_SPI_CCT_N53)
         );
  NAND2XLTF U279 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[0] ), .B(N295), .Y(N32) );
  NAND2XLTF U280 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[1] ), .B(N422), .Y(N35) );
  NAND2XLTF U281 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[3] ), .B(N422), .Y(N41) );
  NAND2XLTF U282 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[4] ), .B(N422), .Y(N44) );
  INVX1TF U283 ( .A(N404), .Y(N407) );
  NAND2XLTF U284 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[2] ), .B(N422), .Y(N38) );
  INVX2TF U285 ( .A(\SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .Y(N367) );
  OAI21XLTF U286 ( .A0(N297), .A1(N285), .B0(N326), .Y(SCPU_CTRL_SPI_CCT_N51)
         );
  NAND2XLTF U287 ( .A(N333), .B(N391), .Y(N332) );
  NAND2XLTF U288 ( .A(SCPU_CTRL_SPI_A_SPI[0]), .B(SCPU_CTRL_SPI_A_SPI[1]), .Y(
        N417) );
  NAND2XLTF U289 ( .A(N102), .B(N284), .Y(N392) );
  NOR2X1TF U290 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .B(
        \SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .Y(N340) );
  CLKBUFX2TF U291 ( .A(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .Y(N390) );
  NOR2X4TF U292 ( .A(SCPU_CTRL_SPI_CEN), .B(N353), .Y(N321) );
  CLKBUFX2TF U293 ( .A(\SCPU_CTRL_SPI_IO_CONTROL[6] ), .Y(N271) );
  INVX2TF U294 ( .A(N390), .Y(N272) );
  INVX2TF U295 ( .A(N390), .Y(N273) );
  NOR3X1TF U296 ( .A(\SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .B(N283), .C(N353), 
        .Y(N324) );
  CLKBUFX2TF U297 ( .A(N241), .Y(N293) );
  INVX2TF U298 ( .A(I_CTRL_BGN), .Y(N274) );
  NOR3X4TF U299 ( .A(N355), .B(N354), .C(N294), .Y(N364) );
  NOR3X2TF U300 ( .A(\SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .B(
        \SCPU_CTRL_SPI_PUT_CNT_STATE[2] ), .C(N288), .Y(N391) );
  INVX2TF U301 ( .A(N426), .Y(N275) );
  NOR2BX1TF U302 ( .AN(N337), .B(N425), .Y(N423) );
  INVX2TF U303 ( .A(I_CTRL_BGN), .Y(N353) );
  NOR2X1TF U304 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ), .B(N298), .Y(N299)
         );
  NAND2X1TF U305 ( .A(N286), .B(N325), .Y(N298) );
  NOR2X1TF U306 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ), .B(N326), .Y(N325)
         );
  NOR2X1TF U307 ( .A(N341), .B(N356), .Y(N352) );
  NAND2X1TF U308 ( .A(N368), .B(I_CTRL_BGN), .Y(N330) );
  NAND2X1TF U309 ( .A(N285), .B(N297), .Y(N326) );
  NAND2X1TF U310 ( .A(N331), .B(N100), .Y(N425) );
  OR2XLTF U311 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[3] ), .B(N271), .Y(N40) );
  OR2XLTF U312 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[0] ), .B(N271), .Y(N31) );
  OR2XLTF U313 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[4] ), .B(N271), .Y(N43) );
  OR2XLTF U314 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[1] ), .B(N271), .Y(N34) );
  OR2XLTF U315 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[2] ), .B(N271), .Y(N37) );
  OAI2BB2XLTF U316 ( .B0(N394), .B1(N393), .A0N(
        \SCPU_CTRL_SPI_PUT_CNT_STATE[2] ), .A1N(N392), .Y(
        SCPU_CTRL_SPI_PUT_N108) );
  NOR2X1TF U317 ( .A(N339), .B(N100), .Y(N354) );
  NOR2X1TF U318 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .B(N280), .Y(N333) );
  NOR2X1TF U319 ( .A(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ), .B(N336), .Y(N341)
         );
  NAND3X1TF U320 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .B(
        \SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .C(N100), .Y(N351) );
  OAI2BB2XLTF U321 ( .B0(N367), .B1(N330), .A0N(N324), .A1N(N323), .Y(N216) );
  NOR2BX1TF U322 ( .AN(N340), .B(N100), .Y(N222) );
  AND2X2TF U323 ( .A(N321), .B(N93), .Y(N322) );
  OAI2BB1X1TF U324 ( .A0N(\SCPU_CTRL_SPI_CCT_REG_BITS[8] ), .A1N(N321), .B0(
        N300), .Y(A_AFTER_MUX[0]) );
  NAND2X1TF U325 ( .A(\SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .B(N283), .Y(N219)
         );
  NAND2X1TF U326 ( .A(N320), .B(N319), .Y(A_AFTER_MUX[8]) );
  NAND2X1TF U327 ( .A(N315), .B(N314), .Y(A_AFTER_MUX[7]) );
  NAND2X1TF U328 ( .A(N313), .B(N312), .Y(A_AFTER_MUX[6]) );
  NAND2X1TF U329 ( .A(N311), .B(N310), .Y(A_AFTER_MUX[5]) );
  NAND2X1TF U330 ( .A(N309), .B(N308), .Y(A_AFTER_MUX[4]) );
  NAND2X1TF U331 ( .A(N307), .B(N306), .Y(A_AFTER_MUX[3]) );
  NAND2X1TF U332 ( .A(N305), .B(N304), .Y(A_AFTER_MUX[2]) );
  NAND2X1TF U333 ( .A(N303), .B(N302), .Y(A_AFTER_MUX[1]) );
  NOR2X2TF U334 ( .A(N380), .B(N301), .Y(N318) );
  NOR2X2TF U335 ( .A(N301), .B(N388), .Y(N316) );
  NAND2X2TF U336 ( .A(SCPU_CTRL_SPI_IS_I_ADDR), .B(N353), .Y(N388) );
  NOR2X2TF U337 ( .A(I_CTRL_BGN), .B(N103), .Y(N317) );
  NAND2X1TF U338 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .B(N280), .Y(N335) );
  NOR2X1TF U339 ( .A(N391), .B(N288), .Y(SCPU_CTRL_SPI_PUT_N106) );
  AOI21X1TF U340 ( .A0(N428), .A1(N279), .B0(N282), .Y(N45) );
  OAI31X1TF U341 ( .A0(N344), .A1(N335), .A2(N337), .B0(N334), .Y(N212) );
  AOI32X1TF U342 ( .A0(N391), .A1(N100), .A2(N333), .B0(N287), .B1(N332), .Y(
        N334) );
  OAI21X1TF U343 ( .A0(N344), .A1(N343), .B0(N342), .Y(N209) );
  OAI21X1TF U344 ( .A0(N287), .A1(N393), .B0(\SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), 
        .Y(N342) );
  AOI211X1TF U345 ( .A0(N341), .A1(N287), .B0(N340), .C0(N275), .Y(N343) );
  AOI22X1TF U346 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .A1(N275), .B0(
        N426), .B1(N281), .Y(N33) );
  OAI32X1TF U347 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ), .A1(
        \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .A2(N426), .B0(N424), .B1(N277), 
        .Y(N36) );
  OAI32X1TF U348 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] ), .A1(N427), .A2(
        N426), .B0(N428), .B1(N279), .Y(N42) );
  NOR2X1TF U349 ( .A(N425), .B(N427), .Y(N428) );
  NOR2X1TF U350 ( .A(N100), .B(N344), .Y(N338) );
  AOI21X1TF U351 ( .A0(N287), .A1(N339), .B0(N391), .Y(N344) );
  NOR2X1TF U352 ( .A(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .B(N425), .Y(N424)
         );
  OAI211X1TF U353 ( .A0(N352), .A1(N290), .B0(N351), .C0(N350), .Y(N205) );
  AOI22X1TF U354 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ), .A1(N346), .B0(
        N347), .B1(N292), .Y(N208) );
  AOI21X1TF U355 ( .A0(N354), .A1(N336), .B0(N394), .Y(N346) );
  OAI211X1TF U356 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .A1(N350), .B0(
        N351), .C0(N349), .Y(N206) );
  OAI21X1TF U357 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .A1(N394), .B0(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .Y(N349) );
  OAI22X1TF U358 ( .A0(I_CTRL_MODE[0]), .A1(N328), .B0(N327), .B1(N330), .Y(
        N215) );
  AOI21X1TF U359 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ), .A1(N326), .B0(
        N325), .Y(N327) );
  OAI21X1TF U360 ( .A0(N383), .A1(N366), .B0(N358), .Y(N202) );
  AOI22X1TF U361 ( .A0(N364), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[2]), .B0(N363), 
        .B1(SCPU_CTRL_SPI_PUT_SRAM_REGS[3]), .Y(N358) );
  OAI21X1TF U362 ( .A0(N381), .A1(N366), .B0(N365), .Y(N197) );
  AOI22X1TF U363 ( .A0(N364), .A1(I_SPI_SO), .B0(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[1]), .B1(N363), .Y(N365) );
  OAI21X1TF U364 ( .A0(N384), .A1(N366), .B0(N359), .Y(N201) );
  AOI22X1TF U365 ( .A0(N364), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[3]), .B0(N363), 
        .B1(SCPU_CTRL_SPI_PUT_SRAM_REGS[4]), .Y(N359) );
  OAI21X1TF U366 ( .A0(N386), .A1(N366), .B0(N361), .Y(N199) );
  AOI22X1TF U367 ( .A0(N364), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[5]), .B0(N363), 
        .B1(SCPU_CTRL_SPI_PUT_SRAM_REGS[6]), .Y(N361) );
  OAI21X1TF U368 ( .A0(N387), .A1(N366), .B0(N362), .Y(N198) );
  AOI22X1TF U369 ( .A0(N364), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[6]), .B0(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[7]), .B1(N363), .Y(N362) );
  OAI21X1TF U370 ( .A0(N382), .A1(N366), .B0(N357), .Y(N203) );
  AOI22X1TF U371 ( .A0(N364), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[1]), .B0(N363), 
        .B1(SCPU_CTRL_SPI_PUT_SRAM_REGS[2]), .Y(N357) );
  OAI21X1TF U372 ( .A0(N385), .A1(N366), .B0(N360), .Y(N200) );
  AOI22X1TF U373 ( .A0(N364), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[4]), .B0(N363), 
        .B1(SCPU_CTRL_SPI_PUT_SRAM_REGS[5]), .Y(N360) );
  NOR2X2TF U374 ( .A(N294), .B(N356), .Y(N363) );
  NAND3X2TF U375 ( .A(N353), .B(N270), .C(N355), .Y(N366) );
  INVX2TF U376 ( .A(N391), .Y(N393) );
  OAI31X1TF U377 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .A1(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .A2(N394), .B0(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ), .Y(N348) );
  NOR2X1TF U378 ( .A(N355), .B(N352), .Y(N394) );
  INVX2TF U379 ( .A(N354), .Y(N356) );
  INVX2TF U380 ( .A(N333), .Y(N339) );
  INVX2TF U381 ( .A(N345), .Y(N336) );
  NOR3X1TF U382 ( .A(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ), .B(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .C(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .Y(N345) );
  INVX2TF U383 ( .A(N351), .Y(N355) );
  INVX2TF U384 ( .A(N330), .Y(N158) );
  OAI21X1TF U385 ( .A0(N381), .A1(N379), .B0(N370), .Y(N196) );
  AOI22X1TF U386 ( .A0(N293), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[1] ), .B0(N377), 
        .B1(I_CTRL_SO), .Y(N370) );
  OAI21X1TF U387 ( .A0(N379), .A1(N384), .B0(N373), .Y(N193) );
  AOI22X1TF U388 ( .A0(N293), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[4] ), .B0(N377), 
        .B1(\SCPU_CTRL_SPI_CCT_REG_BITS[3] ), .Y(N373) );
  OAI21X1TF U389 ( .A0(N379), .A1(N382), .B0(N371), .Y(N195) );
  AOI22X1TF U390 ( .A0(N293), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[2] ), .B0(N377), 
        .B1(\SCPU_CTRL_SPI_CCT_REG_BITS[1] ), .Y(N371) );
  OAI21X1TF U391 ( .A0(N379), .A1(N383), .B0(N372), .Y(N194) );
  AOI22X1TF U392 ( .A0(N293), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[3] ), .B0(N377), 
        .B1(\SCPU_CTRL_SPI_CCT_REG_BITS[2] ), .Y(N372) );
  OAI21X1TF U393 ( .A0(N379), .A1(N385), .B0(N374), .Y(N192) );
  AOI22X1TF U394 ( .A0(N293), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[5] ), .B0(N377), 
        .B1(\SCPU_CTRL_SPI_CCT_REG_BITS[4] ), .Y(N374) );
  OAI21X1TF U395 ( .A0(N379), .A1(N387), .B0(N376), .Y(N190) );
  AOI22X1TF U396 ( .A0(N293), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[7] ), .B0(N377), 
        .B1(\SCPU_CTRL_SPI_CCT_REG_BITS[6] ), .Y(N376) );
  OAI21X1TF U397 ( .A0(N379), .A1(N386), .B0(N375), .Y(N191) );
  AOI22X1TF U398 ( .A0(N293), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[6] ), .B0(N377), 
        .B1(\SCPU_CTRL_SPI_CCT_REG_BITS[5] ), .Y(N375) );
  OAI21X1TF U399 ( .A0(N379), .A1(N389), .B0(N378), .Y(N189) );
  AOI22X1TF U400 ( .A0(N293), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[8] ), .B0(N377), 
        .B1(\SCPU_CTRL_SPI_CCT_REG_BITS[7] ), .Y(N378) );
  NOR2X2TF U401 ( .A(N293), .B(N369), .Y(N377) );
  NAND2X2TF U402 ( .A(I_CTRL_BGN), .B(N369), .Y(N379) );
  NOR3X1TF U403 ( .A(I_CTRL_MODE[1]), .B(N368), .C(N219), .Y(N369) );
  NOR3X1TF U404 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ), .B(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ), .C(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .Y(N297) );
  NOR2X1TF U405 ( .A(N91), .B(\SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .Y(N220) );
  AOI32X1TF U406 ( .A0(N103), .A1(N353), .A2(SCPU_CTRL_SPI_D_WE), .B0(
        I_CTRL_BGN), .B1(N93), .Y(WEN_AFTER_MUX) );
  NOR2X1TF U407 ( .A(N387), .B(N388), .Y(SCPU_CTRL_SPI_I_DATAIN[6]) );
  NOR2X1TF U408 ( .A(N381), .B(N388), .Y(SCPU_CTRL_SPI_I_DATAIN[0]) );
  NOR2X1TF U409 ( .A(N385), .B(N388), .Y(SCPU_CTRL_SPI_I_DATAIN[4]) );
  NOR2X1TF U410 ( .A(N383), .B(N388), .Y(SCPU_CTRL_SPI_I_DATAIN[2]) );
  NOR2X1TF U411 ( .A(N386), .B(N388), .Y(SCPU_CTRL_SPI_I_DATAIN[5]) );
  NOR2X1TF U412 ( .A(N382), .B(N388), .Y(SCPU_CTRL_SPI_I_DATAIN[1]) );
  NOR2X1TF U413 ( .A(N389), .B(N388), .Y(SCPU_CTRL_SPI_I_DATAIN[7]) );
  NOR2X1TF U414 ( .A(N384), .B(N388), .Y(SCPU_CTRL_SPI_I_DATAIN[3]) );
  NOR2X1TF U415 ( .A(N389), .B(N380), .Y(SCPU_CTRL_SPI_D_DATAIN[7]) );
  INVX2TF U416 ( .A(Q_FROM_SRAM[7]), .Y(N389) );
  NOR2X1TF U417 ( .A(N385), .B(N380), .Y(SCPU_CTRL_SPI_D_DATAIN[4]) );
  INVX2TF U418 ( .A(Q_FROM_SRAM[4]), .Y(N385) );
  NOR2X1TF U419 ( .A(N386), .B(N380), .Y(SCPU_CTRL_SPI_D_DATAIN[5]) );
  INVX2TF U420 ( .A(Q_FROM_SRAM[5]), .Y(N386) );
  NOR2X1TF U421 ( .A(N382), .B(N380), .Y(SCPU_CTRL_SPI_D_DATAIN[1]) );
  INVX2TF U422 ( .A(Q_FROM_SRAM[1]), .Y(N382) );
  NOR2X1TF U423 ( .A(N381), .B(N380), .Y(SCPU_CTRL_SPI_D_DATAIN[0]) );
  INVX2TF U424 ( .A(Q_FROM_SRAM[0]), .Y(N381) );
  NOR2X1TF U425 ( .A(N383), .B(N380), .Y(SCPU_CTRL_SPI_D_DATAIN[2]) );
  INVX2TF U426 ( .A(Q_FROM_SRAM[2]), .Y(N383) );
  NOR2X1TF U427 ( .A(N387), .B(N380), .Y(SCPU_CTRL_SPI_D_DATAIN[6]) );
  INVX2TF U428 ( .A(Q_FROM_SRAM[6]), .Y(N387) );
  NOR2X1TF U429 ( .A(N384), .B(N380), .Y(SCPU_CTRL_SPI_D_DATAIN[3]) );
  INVX2TF U430 ( .A(Q_FROM_SRAM[3]), .Y(N384) );
  OAI32X1TF U431 ( .A0(N294), .A1(N331), .A2(N103), .B0(N425), .B1(N294), .Y(
        N213) );
  OAI31X1TF U432 ( .A0(SCPU_CTRL_SPI_A_SPI[1]), .A1(N421), .A2(N291), .B0(N419), .Y(N79) );
  AOI22X1TF U433 ( .A0(SCPU_CTRL_SPI_A_SPI[1]), .A1(N418), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[1] ), .B1(N294), .Y(N419) );
  AOI21X1TF U434 ( .A0(N275), .A1(SCPU_CTRL_SPI_A_SPI[0]), .B0(N295), .Y(N418)
         );
  OAI31X1TF U435 ( .A0(SCPU_CTRL_SPI_A_SPI[3]), .A1(N421), .A2(N414), .B0(N413), .Y(N81) );
  AOI22X1TF U436 ( .A0(SCPU_CTRL_SPI_A_SPI[3]), .A1(N412), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[3] ), .B1(N295), .Y(N413) );
  AOI21X1TF U437 ( .A0(N275), .A1(N411), .B0(N295), .Y(N412) );
  OAI31X1TF U438 ( .A0(SCPU_CTRL_SPI_A_SPI[5]), .A1(N421), .A2(N407), .B0(N406), .Y(N83) );
  AOI22X1TF U439 ( .A0(SCPU_CTRL_SPI_A_SPI[5]), .A1(N405), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[5] ), .B1(N294), .Y(N406) );
  AOI21X1TF U440 ( .A0(N275), .A1(N404), .B0(N295), .Y(N405) );
  OAI31X1TF U441 ( .A0(SCPU_CTRL_SPI_A_SPI[2]), .A1(N421), .A2(N417), .B0(N416), .Y(N80) );
  AOI22X1TF U442 ( .A0(SCPU_CTRL_SPI_A_SPI[2]), .A1(N415), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[2] ), .B1(N295), .Y(N416) );
  AOI31X1TF U443 ( .A0(N275), .A1(SCPU_CTRL_SPI_A_SPI[0]), .A2(
        SCPU_CTRL_SPI_A_SPI[1]), .B0(N295), .Y(N415) );
  OAI31X1TF U444 ( .A0(SCPU_CTRL_SPI_A_SPI[4]), .A1(N421), .A2(N410), .B0(N409), .Y(N82) );
  AOI22X1TF U445 ( .A0(SCPU_CTRL_SPI_A_SPI[4]), .A1(N408), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[4] ), .B1(N295), .Y(N409) );
  AOI31X1TF U446 ( .A0(N275), .A1(N411), .A2(SCPU_CTRL_SPI_A_SPI[3]), .B0(N295), .Y(N408) );
  OAI31X1TF U447 ( .A0(SCPU_CTRL_SPI_A_SPI[6]), .A1(N421), .A2(N403), .B0(N402), .Y(N84) );
  AOI22X1TF U448 ( .A0(SCPU_CTRL_SPI_A_SPI[6]), .A1(N401), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[6] ), .B1(N294), .Y(N402) );
  AOI31X1TF U449 ( .A0(N423), .A1(N404), .A2(SCPU_CTRL_SPI_A_SPI[5]), .B0(N295), .Y(N401) );
  AOI22X1TF U450 ( .A0(N318), .A1(SCPU_CTRL_SPI_D_ADDR[8]), .B0(N321), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[16] ), .Y(N319) );
  AOI22X1TF U451 ( .A0(SCPU_CTRL_SPI_A_SPI[8]), .A1(N317), .B0(N316), .B1(
        SCPU_CTRL_SPI_I_ADDR[8]), .Y(N320) );
  AOI22X1TF U452 ( .A0(N318), .A1(SCPU_CTRL_SPI_D_ADDR[7]), .B0(N321), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[15] ), .Y(N314) );
  AOI22X1TF U453 ( .A0(SCPU_CTRL_SPI_A_SPI[7]), .A1(N317), .B0(N316), .B1(
        SCPU_CTRL_SPI_I_ADDR[7]), .Y(N315) );
  AOI22X1TF U454 ( .A0(N318), .A1(SCPU_CTRL_SPI_D_ADDR[6]), .B0(N321), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[14] ), .Y(N312) );
  AOI22X1TF U455 ( .A0(SCPU_CTRL_SPI_A_SPI[6]), .A1(N317), .B0(N316), .B1(
        SCPU_CTRL_SPI_I_ADDR[6]), .Y(N313) );
  AOI22X1TF U456 ( .A0(N318), .A1(SCPU_CTRL_SPI_D_ADDR[5]), .B0(N321), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[13] ), .Y(N310) );
  AOI22X1TF U457 ( .A0(SCPU_CTRL_SPI_A_SPI[5]), .A1(N317), .B0(N316), .B1(
        SCPU_CTRL_SPI_I_ADDR[5]), .Y(N311) );
  AOI22X1TF U458 ( .A0(N318), .A1(SCPU_CTRL_SPI_D_ADDR[4]), .B0(N321), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[12] ), .Y(N308) );
  AOI22X1TF U459 ( .A0(SCPU_CTRL_SPI_A_SPI[4]), .A1(N317), .B0(N316), .B1(
        SCPU_CTRL_SPI_I_ADDR[4]), .Y(N309) );
  AOI22X1TF U460 ( .A0(N318), .A1(SCPU_CTRL_SPI_D_ADDR[3]), .B0(N321), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[11] ), .Y(N306) );
  AOI22X1TF U461 ( .A0(SCPU_CTRL_SPI_A_SPI[3]), .A1(N317), .B0(N316), .B1(
        SCPU_CTRL_SPI_I_ADDR[3]), .Y(N307) );
  AOI22X1TF U462 ( .A0(N318), .A1(SCPU_CTRL_SPI_D_ADDR[2]), .B0(N321), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[10] ), .Y(N304) );
  AOI22X1TF U463 ( .A0(SCPU_CTRL_SPI_A_SPI[2]), .A1(N317), .B0(N316), .B1(
        SCPU_CTRL_SPI_I_ADDR[2]), .Y(N305) );
  AOI22X1TF U464 ( .A0(N318), .A1(SCPU_CTRL_SPI_D_ADDR[1]), .B0(N321), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[9] ), .Y(N302) );
  AOI22X1TF U465 ( .A0(SCPU_CTRL_SPI_A_SPI[1]), .A1(N317), .B0(N316), .B1(
        SCPU_CTRL_SPI_I_ADDR[1]), .Y(N303) );
  OAI31X1TF U466 ( .A0(SCPU_CTRL_SPI_A_SPI[8]), .A1(N289), .A2(N398), .B0(N397), .Y(N86) );
  AOI22X1TF U467 ( .A0(SCPU_CTRL_SPI_A_SPI[8]), .A1(N396), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[8] ), .B1(N294), .Y(N397) );
  OAI21X1TF U468 ( .A0(SCPU_CTRL_SPI_A_SPI[7]), .A1(N421), .B0(N400), .Y(N396)
         );
  OAI21X1TF U469 ( .A0(N400), .A1(N289), .B0(N399), .Y(N85) );
  INVX2TF U470 ( .A(N414), .Y(N411) );
  OAI21X1TF U471 ( .A0(SCPU_CTRL_SPI_A_SPI[0]), .A1(N421), .B0(N420), .Y(N78)
         );
  INVX2TF U472 ( .A(N423), .Y(N426) );
  NAND2X2TF U473 ( .A(N423), .B(N270), .Y(N421) );
  INVX2TF U474 ( .A(N335), .Y(N331) );
  NOR2X1TF U475 ( .A(N100), .B(N335), .Y(N221) );
  NOR3X1TF U476 ( .A(N102), .B(N103), .C(N284), .Y(I_SCLK1) );
  OAI2BB1X1TF U477 ( .A0N(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .A1N(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ), .B0(N296), .Y(
        SCPU_CTRL_SPI_CCT_N49) );
  OAI221XLTF U478 ( .A0(N103), .A1(SCPU_CTRL_SPI_A_SPI[0]), .B0(N301), .B1(
        SCPU_CTRL_SPI_I_ADDR[0]), .C0(N353), .Y(N300) );
  NOR2BX1TF U479 ( .AN(SCPU_CTRL_SPI_CEN), .B(N353), .Y(CEN_AFTER_MUX) );
  AO22X1TF U480 ( .A0(N322), .A1(I_CTRL_SO), .B0(SCPU_CTRL_SPI_D_DATAOUT[0]), 
        .B1(N353), .Y(D_AFTER_MUX[0]) );
  AO22X1TF U481 ( .A0(N322), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[1] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[1]), .B1(N353), .Y(D_AFTER_MUX[1]) );
  AO22X1TF U482 ( .A0(N322), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[2] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[2]), .B1(N353), .Y(D_AFTER_MUX[2]) );
  AO22X1TF U483 ( .A0(N322), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[3] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[3]), .B1(N274), .Y(D_AFTER_MUX[3]) );
  AO22X1TF U484 ( .A0(N322), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[4] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[4]), .B1(N274), .Y(D_AFTER_MUX[4]) );
  AO22X1TF U485 ( .A0(N322), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[5] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[5]), .B1(N274), .Y(D_AFTER_MUX[5]) );
  AO22X1TF U486 ( .A0(N322), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[6] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[6]), .B1(N274), .Y(D_AFTER_MUX[6]) );
  AO22X1TF U487 ( .A0(N322), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[7] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[7]), .B1(N274), .Y(D_AFTER_MUX[7]) );
  NAND2BX1TF U488 ( .AN(N219), .B(I_CTRL_MODE[1]), .Y(N218) );
  OAI221XLTF U489 ( .A0(\SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .A1(I_LOAD_N), 
        .B0(N367), .B1(N368), .C0(I_CTRL_BGN), .Y(N323) );
  NAND3BX1TF U490 ( .AN(I_LOAD_N), .B(N299), .C(N324), .Y(N328) );
  AO21X1TF U491 ( .A0(I_CTRL_MODE[0]), .A1(I_CTRL_MODE[1]), .B0(N328), .Y(N329) );
  NAND3X1TF U492 ( .A(N278), .B(N281), .C(N277), .Y(N427) );
  NAND3BX1TF U493 ( .AN(N427), .B(N279), .C(N282), .Y(N337) );
  OAI222X1TF U494 ( .A0(N426), .A1(N344), .B0(N339), .B1(N341), .C0(N280), 
        .C1(N338), .Y(N210) );
  NAND2X1TF U495 ( .A(N345), .B(N352), .Y(N347) );
  NAND3X1TF U496 ( .A(N351), .B(N348), .C(N347), .Y(N207) );
  NAND2X1TF U497 ( .A(N352), .B(N290), .Y(N350) );
  OAI2BB2XLTF U498 ( .B0(N389), .B1(N366), .A0N(N364), .A1N(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[7]), .Y(N204) );
  AO22X1TF U499 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[0]), .B0(N273), .B1(I_ADC_PI[0]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[0]) );
  AO22X1TF U500 ( .A0(N390), .A1(SCPU_CTRL_SPI_FOUT[10]), .B0(N272), .B1(
        I_ADC_PI[10]), .Y(SCPU_CTRL_SPI_IO_DATAINA[10]) );
  AO22X1TF U501 ( .A0(N390), .A1(SCPU_CTRL_SPI_FOUT[11]), .B0(N272), .B1(
        I_ADC_PI[11]), .Y(SCPU_CTRL_SPI_IO_DATAINA[11]) );
  AO22X1TF U502 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[12]), .B0(N273), .B1(I_ADC_PI[12]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[12]) );
  NOR2BX1TF U503 ( .AN(I_ADC_PI[13]), .B(N390), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[13]) );
  AO22X1TF U504 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[1]), .B0(N272), .B1(I_ADC_PI[1]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[1]) );
  AO22X1TF U505 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[2]), .B0(N273), .B1(I_ADC_PI[2]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[2]) );
  AO22X1TF U506 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[3]), .B0(N272), .B1(I_ADC_PI[3]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[3]) );
  AO22X1TF U507 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[4]), .B0(N273), .B1(I_ADC_PI[4]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[4]) );
  AO22X1TF U508 ( .A0(N390), .A1(SCPU_CTRL_SPI_FOUT[5]), .B0(N273), .B1(
        I_ADC_PI[5]), .Y(SCPU_CTRL_SPI_IO_DATAINA[5]) );
  AO22X1TF U509 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[6]), .B0(N273), .B1(I_ADC_PI[6]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[6]) );
  AO22X1TF U510 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[7]), .B0(N272), .B1(I_ADC_PI[7]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[7]) );
  AO22X1TF U511 ( .A0(N390), .A1(SCPU_CTRL_SPI_FOUT[8]), .B0(N273), .B1(
        I_ADC_PI[8]), .Y(SCPU_CTRL_SPI_IO_DATAINA[8]) );
  AO22X1TF U512 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[9]), .B0(N273), .B1(I_ADC_PI[9]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[9]) );
  OAI2BB2XLTF U513 ( .B0(N284), .B1(N102), .A0N(N284), .A1N(
        SCPU_CTRL_SPI_PUT_N106), .Y(SCPU_CTRL_SPI_PUT_N107) );
  NAND3X1TF U514 ( .A(SCPU_CTRL_SPI_A_SPI[2]), .B(SCPU_CTRL_SPI_A_SPI[0]), .C(
        SCPU_CTRL_SPI_A_SPI[1]), .Y(N414) );
  NAND2X1TF U515 ( .A(N411), .B(SCPU_CTRL_SPI_A_SPI[3]), .Y(N410) );
  NOR2BX1TF U516 ( .AN(SCPU_CTRL_SPI_A_SPI[4]), .B(N410), .Y(N404) );
  NAND2X1TF U517 ( .A(N404), .B(SCPU_CTRL_SPI_A_SPI[5]), .Y(N403) );
  NOR2BX1TF U518 ( .AN(SCPU_CTRL_SPI_A_SPI[6]), .B(N403), .Y(N395) );
  NAND2BX1TF U519 ( .AN(N421), .B(N395), .Y(N398) );
  OAI2BB1X1TF U520 ( .A0N(N423), .A1N(N395), .B0(N270), .Y(N400) );
  AOI2BB2X1TF U521 ( .B0(\SCPU_CTRL_SPI_IO_DATAOUTA[7] ), .B1(N294), .A0N(
        SCPU_CTRL_SPI_A_SPI[7]), .A1N(N398), .Y(N399) );
endmodule

