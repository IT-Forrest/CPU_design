
module SHARE_SUPERALU_VG ( CLK, RST_N, X_IN, Y_IN, ALU_START, ALU_TYPE, MODE_TYPE, 
        OFFSET, FOUT, POUT, ALU_IS_DONE );
  input [12:0] X_IN;
  input [12:0] Y_IN;
  input [2:0] ALU_TYPE;
  input [1:0] MODE_TYPE;
  input [9:0] OFFSET;
  output [12:0] FOUT;
  output [12:0] POUT;
  input CLK, RST_N, ALU_START;
  output ALU_IS_DONE;
  wire   POST_WORK, PRE_WORK, \INDEX[2] , \RSHT_BITS[3] , SIGN_Y, C152_DATA4_0,
         C152_DATA4_1, C152_DATA4_2, C152_DATA4_3, C152_DATA4_4, C152_DATA4_5,
         C152_DATA4_6, C152_DATA4_7, C152_DATA4_8, C152_DATA4_9, C152_DATA4_10,
         C152_DATA4_11, N73, N74, N90, N91, N92, N121, N122, N123, N124, N128,
         N129, N657, N658, N659, N660, N661, N662, N663, N664, N665, N666,
         N667, N668, N669, N670, N671, N672, N673, N674, N675, N676, N677,
         N678, N679, N680, N681, N682, N683, N684, N685, N686, N687, N688,
         N689, N690, N691, N692, N693, N694, N695, N696, N697, N698, N699,
         N700, N701, N702, N703, N704, N705, N706, N707, N708, N709, N710,
         N711, N712, N713, N714, N715, N716, N717, N718, N719, N720, N721,
         N722, N723, N724, N725, N726, C2_Z_11, C2_Z_10, C2_Z_9, C2_Z_8,
         C2_Z_7, C2_Z_6, C2_Z_5, C2_Z_4, C2_Z_3, C2_Z_2, C2_Z_1, C2_Z_0,
         DP_OP_333_124_4748_N57, DP_OP_333_124_4748_N29,
         DP_OP_333_124_4748_N28, DP_OP_333_124_4748_N27,
         DP_OP_333_124_4748_N26, DP_OP_333_124_4748_N25,
         DP_OP_333_124_4748_N24, DP_OP_333_124_4748_N23,
         DP_OP_333_124_4748_N22, DP_OP_333_124_4748_N21,
         DP_OP_333_124_4748_N20, DP_OP_333_124_4748_N19,
         DP_OP_333_124_4748_N18, DP_OP_333_124_4748_N12,
         DP_OP_333_124_4748_N11, DP_OP_333_124_4748_N10, DP_OP_333_124_4748_N9,
         DP_OP_333_124_4748_N8, DP_OP_333_124_4748_N7, DP_OP_333_124_4748_N6,
         DP_OP_333_124_4748_N5, DP_OP_333_124_4748_N4, DP_OP_333_124_4748_N3,
         DP_OP_333_124_4748_N2, DP_OP_333_124_4748_N1, INTADD_0_CI,
         \INTADD_0_SUM[6] , \INTADD_0_SUM[5] , \INTADD_0_SUM[4] ,
         \INTADD_0_SUM[3] , \INTADD_0_SUM[2] , \INTADD_0_SUM[1] ,
         \INTADD_0_SUM[0] , INTADD_0_N7, INTADD_0_N6, INTADD_0_N5, INTADD_0_N4,
         INTADD_0_N3, INTADD_0_N2, INTADD_0_N1, ADD_X_132_1_N13,
         ADD_X_132_1_N12, ADD_X_132_1_N11, ADD_X_132_1_N10, ADD_X_132_1_N9,
         ADD_X_132_1_N8, ADD_X_132_1_N7, ADD_X_132_1_N6, ADD_X_132_1_N5,
         ADD_X_132_1_N4, ADD_X_132_1_N3, ADD_X_132_1_N2, N1, N2, N3, N4, N5,
         N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N81,
         N82, N83, N84, N85, N86, N87, N88, N89, N93, N94, N95, N96, N97, N98,
         N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N125,
         N126, N127, N130, N131, N132, N133, N134, N135, N136, N137, N138,
         N139, N140, N141, N142, N143, N144, N145, N146, N147, N149, N150,
         N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161,
         N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172,
         N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183,
         N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194,
         N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205,
         N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216,
         N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227,
         N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238,
         N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249,
         N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260,
         N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271,
         N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282,
         N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293,
         N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304,
         N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315,
         N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326,
         N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337,
         N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, N348,
         N349, N350, N351, N352, N353, N354, N355, N356, N357, N358, N359,
         N360, N361, N362, N363, N364, N365, N366, N367, N368, N369, N370,
         N371, N372, N373, N374, N375, N376, N377, N378, N379, N380, N381,
         N382, N383, N384, N385, N386, N387, N388, N389, N390, N391, N392,
         N393, N394, N395, N396, N397, N398, N399, N400, N401, N402, N403,
         N404, N405, N406, N407, N408, N409, N410, N411, N412, N413, N414,
         N415, N416, N417, N418, N419, N420, N421, N422, N423, N424, N425,
         N426, N427, N428, N429, N430, N431, N432, N433, N434, N435, N436,
         N437, N438, N439, N440, N441, N442, N443, N444, N445, N446, N447,
         N448, N449, N450, N451, N452, N453, N454, N455, N456, N457, N458,
         N459, N460, N461, N462, N463, N464, N465, N466, N467, N468, N469,
         N470, N471, N472, N473, N474, N475, N476, N477, N478, N479, N480,
         N481, N482, N483, N484, N485, N486, N487, N488, N489, N490, N491,
         N492, N493, N494, N495, N496, N497, N498, N499, N500, N501, N502,
         N503, N504, N505, N506, N507, N508, N509, N510, N511, N512, N513,
         N514, N515, N516, N517, N518, N519, N520, N521, N522, N523, N524,
         N525, N526, N527, N528, N529, N530, N531, N532, N533, N534, N535,
         N536, N537, N538, N539, N540, N541, N542, N543, N544, N545, N546,
         N547, N548, N549, N550, N551, N552, N553, N554, N555, N556, N557,
         N558, N559, N560, N561, N562, N563, N564, N565, N566, N567, N568,
         N569, N570, N571, N572, N573, N574, N575, N576, N577, N578, N579,
         N580, N581, N582, N583, N584, N585, N586, N587, N588, N589, N590,
         N591, N592, N593, N594, N595, N596, N597, N598, N599, N600, N601,
         N602, N603, N604, N605, N606, N607, N608, N609, N610, N611, N612,
         N613, N614, N615, N616, N617, N618, N619, N620, N621, N622, N623,
         N624, N625, N626, N627, N628, N629, N630, N631, N632, N633, N634,
         N635, N636, N637, N638, N639, N640, N641, N642, N643, N644, N645,
         N646, N647, N648, N649, N650, N651, N652, N653, N654, N655, N656,
         N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737,
         N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748,
         N749, N750, N751, N752, N753, N754, N755, N756, N757, N758, N759,
         N760, N761, N762, N763, N764, N765, N766, N767, N768, N769, N770,
         N771, N772, N773, N774, N775, N776, N777, N778, N779, N780, N781,
         N782, N783, N784, N785, N786, N787, N788, N789, N790, N791, N792,
         N793, N794, N795, N796, N797, N798, N799, N800, N801, N802, N803,
         N804, N805, N806, N807, N808, N809, N810, N811, N812, N813, N814,
         N815, N816, N817, N818, N819, N820, N821, N822, N823, N824, N825,
         N826, N827, N828, N829, N830, N831, N832, N833, N834, N835, N836,
         N837, N838, N839, N840, N841, N842, N843, N844, N845, N846, N847,
         N848, N849, N850, N851, N852, N853, N854, N855, N856, N857, N858,
         N859, N860, N861, N862, N863, N864, N865, N866, N867, N868, N869,
         N870, N871, N872, N873, N874, N875, N876, N877, N878, N879, N880,
         N881, N882, N883, N884, N885, N886, N887, N888, N889, N890, N891,
         N892, N893, N894, N895, N896, N897, N898, N899, N900, N901, N902,
         N903, N904, N905, N906, N907, N908, N909, N910, N911, N912, N913,
         N914, N915, N916, N917, N918, N919, N920, N921, N922, N923, N924,
         N925, N926, N927, N928, N929, N930, N931, N932, N933, N934, N935,
         N936, N937, N938, N939, N940, N941, N942, N943, N944, N945, N946,
         N947, N948, N949, N950, N951, N952, N953, N954, N955, N956, N957,
         N958, N959, N960, N961, N962, N963, N964, N965, N966, N967, N968,
         N969, N970, N971, N972, N973, N974, N975, N976, N977, N978, N979,
         N980, N981, N982, N983, N984, N985, N986, N987, N988, N989, N990,
         N991, N992, N993, N994, N995, N996, N997, N998, N999, N1000, N1001,
         N1002, N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011,
         N1012, N1013, N1014, N1015, N1016, N1017, N1018, N1019;
  wire   [12:9] XTEMP;
  wire   [12:0] DIVISION_HEAD;
  wire   [8:0] DIVISION_REMA;
  wire   [12:0] OPER_A;
  wire   [12:0] OPER_B;
  wire   [12:0] SUM_AB;
  wire   [12:0] ZTEMP;
  wire   [3:2] STEP;

  XOR2X1TF \DP_OP_333_124_4748/U28  ( .A(N81), .B(C2_Z_0), .Y(
        DP_OP_333_124_4748_N29) );
  XOR2X1TF \DP_OP_333_124_4748/U27  ( .A(N81), .B(C2_Z_1), .Y(
        DP_OP_333_124_4748_N28) );
  XOR2X1TF \DP_OP_333_124_4748/U26  ( .A(N81), .B(C2_Z_2), .Y(
        DP_OP_333_124_4748_N27) );
  XOR2X1TF \DP_OP_333_124_4748/U25  ( .A(N971), .B(C2_Z_3), .Y(
        DP_OP_333_124_4748_N26) );
  XOR2X1TF \DP_OP_333_124_4748/U24  ( .A(N81), .B(C2_Z_4), .Y(
        DP_OP_333_124_4748_N25) );
  XOR2X1TF \DP_OP_333_124_4748/U23  ( .A(N81), .B(C2_Z_5), .Y(
        DP_OP_333_124_4748_N24) );
  XOR2X1TF \DP_OP_333_124_4748/U22  ( .A(N81), .B(C2_Z_6), .Y(
        DP_OP_333_124_4748_N23) );
  XOR2X1TF \DP_OP_333_124_4748/U21  ( .A(N971), .B(C2_Z_7), .Y(
        DP_OP_333_124_4748_N22) );
  XOR2X1TF \DP_OP_333_124_4748/U20  ( .A(N81), .B(C2_Z_8), .Y(
        DP_OP_333_124_4748_N21) );
  XOR2X1TF \DP_OP_333_124_4748/U19  ( .A(N971), .B(C2_Z_9), .Y(
        DP_OP_333_124_4748_N20) );
  XOR2X1TF \DP_OP_333_124_4748/U18  ( .A(N81), .B(C2_Z_10), .Y(
        DP_OP_333_124_4748_N19) );
  XOR2X1TF \DP_OP_333_124_4748/U17  ( .A(N971), .B(C2_Z_11), .Y(
        DP_OP_333_124_4748_N18) );
  CMPR32X2TF \DP_OP_333_124_4748/U13  ( .A(DP_OP_333_124_4748_N57), .B(N971), 
        .C(DP_OP_333_124_4748_N29), .CO(DP_OP_333_124_4748_N12), .S(
        C152_DATA4_0) );
  ADDHXLTF \DP_OP_333_124_4748/U12  ( .A(DP_OP_333_124_4748_N28), .B(
        DP_OP_333_124_4748_N12), .CO(DP_OP_333_124_4748_N11), .S(C152_DATA4_1)
         );
  ADDHXLTF \DP_OP_333_124_4748/U11  ( .A(DP_OP_333_124_4748_N27), .B(
        DP_OP_333_124_4748_N11), .CO(DP_OP_333_124_4748_N10), .S(C152_DATA4_2)
         );
  ADDHXLTF \DP_OP_333_124_4748/U10  ( .A(DP_OP_333_124_4748_N26), .B(
        DP_OP_333_124_4748_N10), .CO(DP_OP_333_124_4748_N9), .S(C152_DATA4_3)
         );
  ADDHXLTF \DP_OP_333_124_4748/U9  ( .A(DP_OP_333_124_4748_N25), .B(
        DP_OP_333_124_4748_N9), .CO(DP_OP_333_124_4748_N8), .S(C152_DATA4_4)
         );
  ADDHXLTF \DP_OP_333_124_4748/U8  ( .A(DP_OP_333_124_4748_N24), .B(
        DP_OP_333_124_4748_N8), .CO(DP_OP_333_124_4748_N7), .S(C152_DATA4_5)
         );
  ADDHXLTF \DP_OP_333_124_4748/U7  ( .A(DP_OP_333_124_4748_N23), .B(
        DP_OP_333_124_4748_N7), .CO(DP_OP_333_124_4748_N6), .S(C152_DATA4_6)
         );
  ADDHXLTF \DP_OP_333_124_4748/U6  ( .A(DP_OP_333_124_4748_N22), .B(
        DP_OP_333_124_4748_N6), .CO(DP_OP_333_124_4748_N5), .S(C152_DATA4_7)
         );
  ADDHXLTF \DP_OP_333_124_4748/U5  ( .A(DP_OP_333_124_4748_N21), .B(
        DP_OP_333_124_4748_N5), .CO(DP_OP_333_124_4748_N4), .S(C152_DATA4_8)
         );
  ADDHXLTF \DP_OP_333_124_4748/U4  ( .A(DP_OP_333_124_4748_N20), .B(
        DP_OP_333_124_4748_N4), .CO(DP_OP_333_124_4748_N3), .S(C152_DATA4_9)
         );
  ADDHXLTF \DP_OP_333_124_4748/U3  ( .A(DP_OP_333_124_4748_N19), .B(
        DP_OP_333_124_4748_N3), .CO(DP_OP_333_124_4748_N2), .S(C152_DATA4_10)
         );
  ADDHXLTF \DP_OP_333_124_4748/U2  ( .A(DP_OP_333_124_4748_N18), .B(
        DP_OP_333_124_4748_N2), .CO(DP_OP_333_124_4748_N1), .S(C152_DATA4_11)
         );
  CMPR32X2TF \intadd_0/U8  ( .A(X_IN[1]), .B(DIVISION_HEAD[5]), .C(INTADD_0_CI), .CO(INTADD_0_N7), .S(\INTADD_0_SUM[0] ) );
  CMPR32X2TF \intadd_0/U7  ( .A(X_IN[2]), .B(DIVISION_HEAD[6]), .C(INTADD_0_N7), .CO(INTADD_0_N6), .S(\INTADD_0_SUM[1] ) );
  CMPR32X2TF \intadd_0/U6  ( .A(N94), .B(DIVISION_HEAD[7]), .C(INTADD_0_N6), 
        .CO(INTADD_0_N5), .S(\INTADD_0_SUM[2] ) );
  CMPR32X2TF \intadd_0/U5  ( .A(X_IN[4]), .B(DIVISION_HEAD[8]), .C(INTADD_0_N5), .CO(INTADD_0_N4), .S(\INTADD_0_SUM[3] ) );
  CMPR32X2TF \intadd_0/U4  ( .A(N106), .B(DIVISION_HEAD[9]), .C(INTADD_0_N4), 
        .CO(INTADD_0_N3), .S(\INTADD_0_SUM[4] ) );
  CMPR32X2TF \intadd_0/U3  ( .A(X_IN[6]), .B(DIVISION_HEAD[10]), .C(
        INTADD_0_N3), .CO(INTADD_0_N2), .S(\INTADD_0_SUM[5] ) );
  CMPR32X2TF \intadd_0/U2  ( .A(X_IN[7]), .B(DIVISION_HEAD[11]), .C(
        INTADD_0_N2), .CO(INTADD_0_N1), .S(\INTADD_0_SUM[6] ) );
  DFFRX2TF \rsht_bits_reg[3]  ( .D(N704), .CK(CLK), .RN(RST_N), .Q(
        \RSHT_BITS[3] ), .QN(N194) );
  DFFRX2TF \wtemp_reg[9]  ( .D(N673), .CK(CLK), .RN(RST_N), .Q(OPER_B[9]), 
        .QN(N193) );
  DFFRX2TF \wtemp_reg[12]  ( .D(N724), .CK(CLK), .RN(RST_N), .Q(OPER_B[12]), 
        .QN(N192) );
  DFFRX2TF \index_reg[3]  ( .D(N725), .CK(CLK), .RN(RST_N), .Q(N191), .QN(N124) );
  DFFRX2TF \wtemp_reg[11]  ( .D(N671), .CK(CLK), .RN(RST_N), .Q(OPER_B[11]), 
        .QN(N190) );
  DFFRX2TF \wtemp_reg[0]  ( .D(N682), .CK(CLK), .RN(RST_N), .Q(OPER_B[0]), 
        .QN(N189) );
  DFFRX2TF \wtemp_reg[3]  ( .D(N679), .CK(CLK), .RN(RST_N), .Q(OPER_B[3]), 
        .QN(N188) );
  DFFRX2TF \wtemp_reg[1]  ( .D(N681), .CK(CLK), .RN(RST_N), .Q(OPER_B[1]), 
        .QN(N187) );
  DFFRX2TF \index_reg[1]  ( .D(N699), .CK(CLK), .RN(RST_N), .Q(N186), .QN(N128) );
  DFFRX2TF \rsht_bits_reg[0]  ( .D(N703), .CK(CLK), .RN(RST_N), .Q(N185), .QN(
        N92) );
  DFFRX2TF \ytemp_reg[1]  ( .D(N693), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[1]), .QN(N184) );
  DFFRX2TF \ytemp_reg[0]  ( .D(N705), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[0]), .QN(N183) );
  DFFRX2TF sign_y_reg ( .D(N694), .CK(CLK), .RN(RST_N), .Q(SIGN_Y), .QN(N182)
         );
  DFFRX2TF \wtemp_reg[4]  ( .D(N678), .CK(CLK), .RN(RST_N), .Q(OPER_B[4]), 
        .QN(N181) );
  DFFSX2TF pre_work_reg ( .D(N695), .CK(CLK), .SN(RST_N), .Q(PRE_WORK), .QN(
        N180) );
  DFFRX2TF \xtemp_reg[12]  ( .D(N723), .CK(CLK), .RN(RST_N), .Q(XTEMP[12]), 
        .QN(N179) );
  DFFRX2TF \xtemp_reg[8]  ( .D(N711), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[12]), .QN(N178) );
  DFFRX2TF \ytemp_reg[6]  ( .D(N688), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[6]), .QN(N177) );
  DFFRX2TF \ytemp_reg[4]  ( .D(N690), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[4]), .QN(N176) );
  DFFRX2TF \ytemp_reg[10]  ( .D(N684), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[1]), .QN(N175) );
  DFFRX2TF \ytemp_reg[9]  ( .D(N685), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[0]), .QN(N174) );
  DFFRX2TF \ytemp_reg[7]  ( .D(N687), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[7]), .QN(N173) );
  DFFRX2TF \ytemp_reg[5]  ( .D(N689), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[5]), .QN(N172) );
  DFFRX2TF \ytemp_reg[3]  ( .D(N691), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[3]), .QN(N171) );
  DFFRX2TF \step_reg[0]  ( .D(N697), .CK(CLK), .RN(RST_N), .Q(N170), .QN(N122)
         );
  DFFRX2TF \ytemp_reg[11]  ( .D(N683), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[2]), .QN(N168) );
  DFFRX2TF SEL_SRC_reg ( .D(N720), .CK(CLK), .RN(RST_N), .Q(POST_WORK), .QN(
        N167) );
  DFFRX2TF \wtemp_reg[10]  ( .D(N672), .CK(CLK), .RN(RST_N), .Q(OPER_B[10]), 
        .QN(N166) );
  DFFRX2TF \wtemp_reg[8]  ( .D(N674), .CK(CLK), .RN(RST_N), .Q(OPER_B[8]), 
        .QN(N165) );
  DFFRX2TF \rsht_bits_reg[1]  ( .D(N702), .CK(CLK), .RN(RST_N), .Q(N164), .QN(
        N91) );
  DFFRX2TF \index_reg[0]  ( .D(N726), .CK(CLK), .RN(RST_N), .Q(N163), .QN(N129) );
  DFFRX2TF \wtemp_reg[2]  ( .D(N680), .CK(CLK), .RN(RST_N), .Q(OPER_B[2]), 
        .QN(N162) );
  DFFRX2TF \xtemp_reg[10]  ( .D(N709), .CK(CLK), .RN(RST_N), .Q(XTEMP[10]), 
        .QN(N161) );
  DFFRX2TF \xtemp_reg[6]  ( .D(N713), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[10]), .QN(N160) );
  DFFRX2TF \xtemp_reg[11]  ( .D(N708), .CK(CLK), .RN(RST_N), .Q(XTEMP[11]), 
        .QN(N159) );
  DFFRX2TF \xtemp_reg[0]  ( .D(N719), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[4]), .QN(N158) );
  DFFRX2TF \xtemp_reg[2]  ( .D(N717), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[6]), .QN(N157) );
  DFFRX2TF \xtemp_reg[5]  ( .D(N714), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[9]), .QN(N156) );
  DFFRX2TF \xtemp_reg[4]  ( .D(N715), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[8]), .QN(N155) );
  DFFRX2TF \xtemp_reg[7]  ( .D(N712), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[11]), .QN(N154) );
  DFFRX2TF XOR_SRC_reg ( .D(N707), .CK(CLK), .RN(RST_N), .Q(N61), .QN(N73) );
  DFFRX2TF \step_reg[3]  ( .D(N721), .CK(CLK), .RN(RST_N), .Q(STEP[3]), .QN(
        N153) );
  DFFRX2TF \step_reg[1]  ( .D(N700), .CK(CLK), .RN(RST_N), .Q(N152), .QN(N121)
         );
  DFFRX2TF \step_reg[2]  ( .D(N696), .CK(CLK), .RN(RST_N), .Q(STEP[2]), .QN(
        N151) );
  DFFRX2TF \ytemp_reg[2]  ( .D(N692), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[2]), .QN(N150) );
  DFFRX2TF \ytemp_reg[8]  ( .D(N686), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[8]), .QN(N149) );
  DFFRX2TF \rsht_bits_reg[2]  ( .D(N701), .CK(CLK), .RN(RST_N), .QN(N90) );
  DFFRX2TF SEL_Z_reg ( .D(N670), .CK(CLK), .RN(RST_N), .Q(N169), .QN(N123) );
  CMPR32X2TF \add_x_132_1/U4  ( .A(OPER_A[10]), .B(OPER_B[10]), .C(
        ADD_X_132_1_N4), .CO(ADD_X_132_1_N3), .S(SUM_AB[10]) );
  CMPR32X2TF \add_x_132_1/U6  ( .A(OPER_A[8]), .B(OPER_B[8]), .C(
        ADD_X_132_1_N6), .CO(ADD_X_132_1_N5), .S(SUM_AB[8]) );
  CMPR32X2TF \add_x_132_1/U8  ( .A(OPER_A[6]), .B(OPER_B[6]), .C(
        ADD_X_132_1_N8), .CO(ADD_X_132_1_N7), .S(SUM_AB[6]) );
  CMPR32X2TF \add_x_132_1/U10  ( .A(OPER_A[4]), .B(OPER_B[4]), .C(
        ADD_X_132_1_N10), .CO(ADD_X_132_1_N9), .S(SUM_AB[4]) );
  CMPR32X2TF \add_x_132_1/U13  ( .A(OPER_A[1]), .B(OPER_B[1]), .C(
        ADD_X_132_1_N13), .CO(ADD_X_132_1_N12), .S(SUM_AB[1]) );
  CMPR32X2TF \add_x_132_1/U5  ( .A(OPER_A[9]), .B(OPER_B[9]), .C(
        ADD_X_132_1_N5), .CO(ADD_X_132_1_N4), .S(SUM_AB[9]) );
  CMPR32X2TF \add_x_132_1/U12  ( .A(OPER_A[2]), .B(OPER_B[2]), .C(
        ADD_X_132_1_N12), .CO(ADD_X_132_1_N11), .S(SUM_AB[2]) );
  CMPR32X2TF \add_x_132_1/U11  ( .A(OPER_A[3]), .B(OPER_B[3]), .C(
        ADD_X_132_1_N11), .CO(ADD_X_132_1_N10), .S(SUM_AB[3]) );
  CMPR32X2TF \add_x_132_1/U9  ( .A(OPER_A[5]), .B(OPER_B[5]), .C(
        ADD_X_132_1_N9), .CO(ADD_X_132_1_N8), .S(SUM_AB[5]) );
  CMPR32X2TF \add_x_132_1/U7  ( .A(OPER_A[7]), .B(OPER_B[7]), .C(
        ADD_X_132_1_N7), .CO(ADD_X_132_1_N6), .S(SUM_AB[7]) );
  CMPR32X2TF \add_x_132_1/U3  ( .A(OPER_A[11]), .B(OPER_B[11]), .C(
        ADD_X_132_1_N3), .CO(ADD_X_132_1_N2), .S(SUM_AB[11]) );
  DFFRX2TF sign_x_reg ( .D(N722), .CK(CLK), .RN(RST_N), .Q(N965), .QN(N74) );
  DFFRX1TF \wtemp_reg[6]  ( .D(N676), .CK(CLK), .RN(RST_N), .Q(OPER_B[6]) );
  DFFRX1TF \ztemp_reg[0]  ( .D(N669), .CK(CLK), .RN(RST_N), .Q(ZTEMP[0]) );
  DFFRX1TF \ztemp_reg[6]  ( .D(N663), .CK(CLK), .RN(RST_N), .Q(ZTEMP[6]) );
  DFFRX1TF \ztemp_reg[4]  ( .D(N665), .CK(CLK), .RN(RST_N), .Q(ZTEMP[4]) );
  DFFRX1TF \ztemp_reg[2]  ( .D(N667), .CK(CLK), .RN(RST_N), .Q(ZTEMP[2]) );
  DFFRX1TF \ztemp_reg[1]  ( .D(N668), .CK(CLK), .RN(RST_N), .Q(ZTEMP[1]) );
  DFFRX1TF \ztemp_reg[5]  ( .D(N664), .CK(CLK), .RN(RST_N), .Q(ZTEMP[5]) );
  DFFRX1TF \ztemp_reg[3]  ( .D(N666), .CK(CLK), .RN(RST_N), .Q(ZTEMP[3]) );
  DFFRX1TF \ztemp_reg[7]  ( .D(N662), .CK(CLK), .RN(RST_N), .Q(ZTEMP[7]) );
  DFFRX1TF \ztemp_reg[8]  ( .D(N661), .CK(CLK), .RN(RST_N), .Q(ZTEMP[8]) );
  DFFRX1TF \ztemp_reg[9]  ( .D(N660), .CK(CLK), .RN(RST_N), .Q(ZTEMP[9]) );
  DFFRX1TF \wtemp_reg[5]  ( .D(N677), .CK(CLK), .RN(RST_N), .Q(OPER_B[5]) );
  DFFRX1TF \wtemp_reg[7]  ( .D(N675), .CK(CLK), .RN(RST_N), .Q(OPER_B[7]) );
  DFFRX1TF \ztemp_reg[10]  ( .D(N659), .CK(CLK), .RN(RST_N), .Q(ZTEMP[10]) );
  DFFRX1TF \ztemp_reg[11]  ( .D(N658), .CK(CLK), .RN(RST_N), .Q(ZTEMP[11]) );
  DFFRX1TF \ztemp_reg[12]  ( .D(N657), .CK(CLK), .RN(RST_N), .Q(ZTEMP[12]) );
  DFFRX1TF \ytemp_reg[12]  ( .D(N706), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[3]), .QN(N649) );
  DFFRX2TF \xtemp_reg[1]  ( .D(N718), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[5]), .QN(N514) );
  DFFRX2TF \xtemp_reg[9]  ( .D(N710), .CK(CLK), .RN(RST_N), .Q(XTEMP[9]), .QN(
        N529) );
  DFFRX2TF \xtemp_reg[3]  ( .D(N716), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[7]), .QN(N423) );
  DFFRX2TF \index_reg[2]  ( .D(N698), .CK(CLK), .RN(RST_N), .Q(\INDEX[2] ) );
  NAND2X1TF U3 ( .A(N774), .B(N766), .Y(N394) );
  NAND2X1TF U4 ( .A(ALU_START), .B(N263), .Y(N600) );
  OAI21X1TF U5 ( .A0(N893), .A1(N934), .B0(N932), .Y(N1) );
  AO21X1TF U6 ( .A0(N892), .A1(N937), .B0(N890), .Y(N2) );
  AOI22X1TF U7 ( .A0(OPER_A[7]), .A1(N1), .B0(OPER_B[7]), .B1(N2), .Y(N3) );
  OAI31X1TF U8 ( .A0(N892), .A1(N115), .A2(OPER_B[7]), .B0(N3), .Y(N4) );
  AOI211X1TF U9 ( .A0(C152_DATA4_7), .A1(N113), .B0(N211), .C0(N4), .Y(N5) );
  NAND3BX1TF U10 ( .AN(OPER_A[7]), .B(N893), .C(N931), .Y(N6) );
  OAI211X1TF U11 ( .A0(N894), .A1(N165), .B0(N5), .C0(N6), .Y(N675) );
  OAI211X1TF U12 ( .A0(N823), .A1(N376), .B0(N612), .C0(N640), .Y(N7) );
  AOI21XLTF U13 ( .A0(N377), .A1(N822), .B0(N7), .Y(N8) );
  NAND3X1TF U14 ( .A(N378), .B(N543), .C(N8), .Y(N9) );
  OAI22X1TF U15 ( .A0(N640), .A1(N764), .B0(N119), .B1(N379), .Y(N10) );
  OAI21X1TF U16 ( .A0(N10), .A1(N747), .B0(N9), .Y(N11) );
  OAI21X1TF U17 ( .A0(N167), .A1(N9), .B0(N11), .Y(N720) );
  AOI32X1TF U18 ( .A0(N116), .A1(N843), .A2(N935), .B0(N189), .B1(N843), .Y(
        N12) );
  AOI211X1TF U19 ( .A0(C152_DATA4_0), .A1(N114), .B0(N891), .C0(N12), .Y(N13)
         );
  OAI21X1TF U20 ( .A0(N854), .A1(N931), .B0(OPER_A[0]), .Y(N14) );
  OAI211X1TF U21 ( .A0(N187), .A1(N894), .B0(N13), .C0(N14), .Y(N682) );
  AOI22X1TF U22 ( .A0(N1011), .A1(ZTEMP[0]), .B0(N107), .B1(DIVISION_HEAD[0]), 
        .Y(N15) );
  AOI32XLTF U23 ( .A0(N1010), .A1(N15), .A2(N1019), .B0(N976), .B1(N15), .Y(
        N669) );
  OAI32X1TF U24 ( .A0(N190), .A1(N936), .A2(N116), .B0(N935), .B1(N190), .Y(
        N16) );
  CLKINVX1TF U25 ( .A(OPER_A[11]), .Y(N17) );
  OAI32X1TF U26 ( .A0(N17), .A1(N934), .A2(N933), .B0(N932), .B1(N17), .Y(N18)
         );
  AOI31X1TF U27 ( .A0(N933), .A1(N931), .A2(N17), .B0(N930), .Y(N19) );
  NOR2X1TF U28 ( .A(N115), .B(OPER_B[11]), .Y(N20) );
  AOI222XLTF U29 ( .A0(C152_DATA4_11), .A1(N113), .B0(N225), .B1(N964), .C0(
        N936), .C1(N20), .Y(N21) );
  OAI211X1TF U30 ( .A0(N192), .A1(N938), .B0(N19), .C0(N21), .Y(N22) );
  OR3X1TF U31 ( .A(N16), .B(N18), .C(N22), .Y(N671) );
  NOR2X1TF U32 ( .A(N933), .B(OPER_A[11]), .Y(N23) );
  XNOR2X1TF U33 ( .A(OPER_A[12]), .B(N23), .Y(N24) );
  AOI22X1TF U34 ( .A0(N24), .A1(N931), .B0(OPER_A[12]), .B1(N854), .Y(N25) );
  OAI21X1TF U35 ( .A0(N132), .A1(N549), .B0(N140), .Y(N26) );
  XNOR2X1TF U36 ( .A(N26), .B(N971), .Y(N27) );
  XNOR2X1TF U37 ( .A(DP_OP_333_124_4748_N1), .B(N27), .Y(N28) );
  NOR2X1TF U38 ( .A(OPER_B[11]), .B(N936), .Y(N29) );
  OAI31X1TF U39 ( .A0(N115), .A1(N29), .A2(OPER_B[12]), .B0(N825), .Y(N30) );
  AOI211X1TF U40 ( .A0(N114), .A1(N28), .B0(N930), .C0(N30), .Y(N31) );
  OAI31X1TF U41 ( .A0(OPER_B[11]), .A1(N936), .A2(N911), .B0(N874), .Y(N32) );
  AOI32X1TF U42 ( .A0(N130), .A1(OPER_B[12]), .A2(N32), .B0(N222), .B1(
        OPER_B[12]), .Y(N33) );
  NAND4BX1TF U43 ( .AN(N821), .B(N25), .C(N31), .D(N33), .Y(N724) );
  NOR3X1TF U44 ( .A(Y_IN[12]), .B(Y_IN[11]), .C(Y_IN[10]), .Y(N34) );
  NOR2X1TF U45 ( .A(N502), .B(N89), .Y(N35) );
  CLKINVX1TF U46 ( .A(Y_IN[6]), .Y(N36) );
  CLKINVX1TF U47 ( .A(N442), .Y(N37) );
  AOI22X1TF U48 ( .A0(N318), .A1(N37), .B0(N105), .B1(N738), .Y(N38) );
  OAI21X1TF U49 ( .A0(X_IN[4]), .A1(N317), .B0(N93), .Y(N39) );
  OAI22X1TF U50 ( .A0(N105), .A1(N738), .B0(X_IN[6]), .B1(N731), .Y(N40) );
  AOI31X1TF U51 ( .A0(N319), .A1(N38), .A2(N39), .B0(N40), .Y(N41) );
  AOI21X1TF U52 ( .A0(N731), .A1(X_IN[6]), .B0(N41), .Y(N42) );
  OA22X1TF U53 ( .A0(N43), .A1(N42), .B0(N488), .B1(N197), .Y(N44) );
  AO21X1TF U54 ( .A0(N468), .A1(N42), .B0(Y_IN[4]), .Y(N45) );
  AOI22X1TF U55 ( .A0(N488), .A1(N197), .B0(N44), .B1(N45), .Y(N46) );
  OA21XLTF U56 ( .A0(N36), .A1(N46), .B0(X_IN[9]), .Y(N47) );
  AOI211X1TF U57 ( .A0(N46), .A1(N36), .B0(N47), .C0(N35), .Y(N48) );
  AOI21X1TF U58 ( .A0(N502), .A1(Y_IN[7]), .B0(N48), .Y(N49) );
  AOI222XLTF U59 ( .A0(N762), .A1(N138), .B0(N762), .B1(N49), .C0(N138), .C1(
        N49), .Y(N50) );
  OAI21X1TF U60 ( .A0(Y_IN[9]), .A1(N305), .B0(N50), .Y(N51) );
  OAI211X1TF U61 ( .A0(X_IN[12]), .A1(N784), .B0(N34), .C0(N51), .Y(N770) );
  CLKINVX1TF U62 ( .A(X_IN[7]), .Y(N43) );
  NOR3X1TF U63 ( .A(N910), .B(N74), .C(N907), .Y(N52) );
  NOR2X1TF U64 ( .A(N166), .B(N938), .Y(N53) );
  AOI211X1TF U65 ( .A0(N113), .A1(C152_DATA4_9), .B0(N52), .C0(N53), .Y(N54)
         );
  NOR2X1TF U66 ( .A(N934), .B(OPER_A[9]), .Y(N55) );
  AOI22X1TF U67 ( .A0(SIGN_Y), .A1(N906), .B0(N909), .B1(N55), .Y(N56) );
  OAI21X1TF U68 ( .A0(N116), .A1(N908), .B0(N935), .Y(N57) );
  OAI21X1TF U69 ( .A0(N934), .A1(N909), .B0(N932), .Y(N58) );
  AOI22X1TF U70 ( .A0(OPER_B[9]), .A1(N57), .B0(OPER_A[9]), .B1(N58), .Y(N59)
         );
  NAND3X1TF U71 ( .A(N937), .B(N908), .C(N193), .Y(N60) );
  NAND4X1TF U72 ( .A(N54), .B(N56), .C(N59), .D(N60), .Y(N673) );
  INVX2TF U73 ( .A(N941), .Y(N118) );
  NOR3BX2TF U74 ( .AN(ALU_TYPE[2]), .B(ALU_TYPE[0]), .C(ALU_TYPE[1]), .Y(N263)
         );
  NOR3BXLTF U75 ( .AN(ALU_TYPE[0]), .B(ALU_TYPE[1]), .C(ALU_TYPE[2]), .Y(N262)
         );
  OAI32X4TF U76 ( .A0(N768), .A1(N767), .A2(X_IN[0]), .B0(N766), .B1(N768), 
        .Y(N771) );
  NOR2X4TF U77 ( .A(N385), .B(N769), .Y(N807) );
  NAND2X2TF U78 ( .A(PRE_WORK), .B(N971), .Y(N385) );
  OA21XLTF U79 ( .A0(SUM_AB[12]), .A1(N651), .B0(N119), .Y(N144) );
  NAND2X1TF U80 ( .A(N929), .B(N208), .Y(N221) );
  CLKINVX1TF U81 ( .A(SUM_AB[4]), .Y(N388) );
  AO21X1TF U82 ( .A0(N777), .A1(N376), .B0(N823), .Y(N509) );
  CLKAND2X2TF U83 ( .A(N647), .B(N640), .Y(N546) );
  CLKINVX1TF U84 ( .A(N867), .Y(N865) );
  OR3X1TF U85 ( .A(PRE_WORK), .B(N606), .C(N600), .Y(N501) );
  CLKINVX1TF U86 ( .A(Y_IN[6]), .Y(N204) );
  AND2X2TF U87 ( .A(N117), .B(N195), .Y(N245) );
  AND2X2TF U88 ( .A(N195), .B(N73), .Y(N244) );
  CLKINVX1TF U89 ( .A(N839), .Y(N834) );
  CLKINVX1TF U90 ( .A(N197), .Y(N205) );
  CLKINVX1TF U91 ( .A(N621), .Y(N623) );
  AOI211X1TF U92 ( .A0(N94), .A1(N747), .B0(N440), .C0(N439), .Y(N441) );
  AOI211X1TF U93 ( .A0(N106), .A1(N747), .B0(N458), .C0(N457), .Y(N459) );
  AOI211X1TF U94 ( .A0(N89), .A1(N747), .B0(N788), .C0(N787), .Y(N789) );
  OA21XLTF U95 ( .A0(SUM_AB[12]), .A1(N393), .B0(N119), .Y(N505) );
  CLKINVX2TF U96 ( .A(N871), .Y(N215) );
  AOI21X1TF U97 ( .A0(N767), .A1(N309), .B0(N385), .Y(N381) );
  AND2X2TF U98 ( .A(N904), .B(N922), .Y(N937) );
  INVX1TF U99 ( .A(N906), .Y(N889) );
  OR2X2TF U100 ( .A(N1011), .B(N133), .Y(N1012) );
  OAI21XLTF U101 ( .A0(N312), .A1(N629), .B0(N622), .Y(N313) );
  AOI22X1TF U102 ( .A0(Y_IN[9]), .A1(N802), .B0(X_IN[4]), .B1(N136), .Y(N803)
         );
  AOI21X1TF U103 ( .A0(N643), .A1(N130), .B0(N642), .Y(N646) );
  AOI211X2TF U104 ( .A0(N571), .A1(N130), .B0(N595), .C0(N570), .Y(N597) );
  INVX1TF U105 ( .A(N403), .Y(N404) );
  NAND3XLTF U106 ( .A(N130), .B(N824), .C(N823), .Y(N633) );
  OAI31XLTF U107 ( .A0(N119), .A1(N170), .A2(N632), .B0(N631), .Y(N637) );
  OR2X2TF U108 ( .A(N385), .B(N764), .Y(N801) );
  OAI31X1TF U109 ( .A0(N565), .A1(N566), .A2(N564), .B0(N130), .Y(N582) );
  AOI32XLTF U110 ( .A0(N822), .A1(N130), .A2(N823), .B0(N638), .B1(N130), .Y(
        N644) );
  NAND4XLTF U111 ( .A(N612), .B(N611), .C(N610), .D(N609), .Y(N613) );
  OAI2BB2XLTF U112 ( .B0(N762), .B1(N804), .A0N(Y_IN[6]), .A1N(N802), .Y(N779)
         );
  AOI22X1TF U113 ( .A0(X_IN[2]), .A1(N802), .B0(N94), .B1(N444), .Y(N425) );
  AOI22X1TF U114 ( .A0(XTEMP[10]), .A1(N95), .B0(X_IN[7]), .B1(N802), .Y(N480)
         );
  AOI22X1TF U115 ( .A0(X_IN[2]), .A1(N444), .B0(X_IN[1]), .B1(N802), .Y(N417)
         );
  INVX1TF U116 ( .A(OPER_A[10]), .Y(N915) );
  OAI211XLTF U117 ( .A0(N132), .A1(N368), .B0(N973), .C0(N601), .Y(N370) );
  NAND3BXLTF U118 ( .AN(N380), .B(N777), .C(N639), .Y(N369) );
  AOI22X1TF U119 ( .A0(N197), .A1(N802), .B0(N89), .B1(N791), .Y(N755) );
  AOI22X1TF U120 ( .A0(Y_IN[1]), .A1(N802), .B0(DIVISION_REMA[4]), .B1(N125), 
        .Y(N732) );
  INVX1TF U121 ( .A(OPER_A[8]), .Y(N897) );
  INVX2TF U122 ( .A(N736), .Y(N97) );
  INVX1TF U123 ( .A(OPER_A[6]), .Y(N881) );
  INVX1TF U124 ( .A(OPER_A[4]), .Y(N862) );
  AOI22X1TF U125 ( .A0(Y_IN[3]), .A1(N802), .B0(DIVISION_REMA[6]), .B1(N125), 
        .Y(N742) );
  CLKINVX1TF U126 ( .A(OPER_A[1]), .Y(N832) );
  AOI22X1TF U127 ( .A0(DIVISION_HEAD[2]), .A1(N125), .B0(Y_IN[8]), .B1(N802), 
        .Y(N795) );
  INVX2TF U128 ( .A(N132), .Y(N81) );
  INVX2TF U129 ( .A(N747), .Y(N99) );
  AOI22X1TF U130 ( .A0(DIVISION_HEAD[3]), .A1(N110), .B0(ZTEMP[12]), .B1(N143), 
        .Y(N260) );
  AND2X2TF U131 ( .A(N382), .B(N354), .Y(N736) );
  AOI22X1TF U132 ( .A0(DIVISION_HEAD[2]), .A1(N110), .B0(ZTEMP[11]), .B1(N143), 
        .Y(N258) );
  AOI22X1TF U133 ( .A0(DIVISION_HEAD[1]), .A1(N110), .B0(ZTEMP[10]), .B1(N143), 
        .Y(N257) );
  AOI22X1TF U134 ( .A0(DIVISION_HEAD[0]), .A1(N110), .B0(ZTEMP[9]), .B1(N143), 
        .Y(N256) );
  AOI22X1TF U135 ( .A0(DIVISION_REMA[8]), .A1(N110), .B0(ZTEMP[8]), .B1(N169), 
        .Y(N255) );
  AOI22X1TF U136 ( .A0(DIVISION_REMA[7]), .A1(N110), .B0(ZTEMP[7]), .B1(N169), 
        .Y(N254) );
  AOI22X1TF U137 ( .A0(DIVISION_REMA[6]), .A1(N110), .B0(ZTEMP[6]), .B1(N169), 
        .Y(N253) );
  AOI22X1TF U138 ( .A0(DIVISION_REMA[5]), .A1(N110), .B0(ZTEMP[5]), .B1(N169), 
        .Y(N252) );
  AOI22X1TF U139 ( .A0(DIVISION_REMA[4]), .A1(N110), .B0(ZTEMP[4]), .B1(N169), 
        .Y(N251) );
  AOI22X1TF U140 ( .A0(DIVISION_REMA[3]), .A1(N110), .B0(ZTEMP[3]), .B1(N169), 
        .Y(N250) );
  AOI22X1TF U141 ( .A0(DIVISION_REMA[2]), .A1(N109), .B0(ZTEMP[2]), .B1(N169), 
        .Y(N249) );
  AOI22X1TF U142 ( .A0(DIVISION_REMA[1]), .A1(N109), .B0(ZTEMP[1]), .B1(N169), 
        .Y(N248) );
  AOI22X1TF U143 ( .A0(DIVISION_REMA[0]), .A1(N109), .B0(ZTEMP[0]), .B1(N169), 
        .Y(N247) );
  OAI21XLTF U144 ( .A0(N132), .A1(N727), .B0(N207), .Y(C2_Z_0) );
  INVX2TF U145 ( .A(N813), .Y(N120) );
  INVX2TF U146 ( .A(N259), .Y(N109) );
  OAI22X1TF U147 ( .A0(N133), .A1(N805), .B0(OFFSET[9]), .B1(N140), .Y(C2_Z_11) );
  OAI22X1TF U148 ( .A0(N133), .A1(N762), .B0(OFFSET[6]), .B1(N207), .Y(C2_Z_8)
         );
  OAI22X1TF U149 ( .A0(N133), .A1(N784), .B0(OFFSET[7]), .B1(N207), .Y(C2_Z_9)
         );
  OAI22X1TF U150 ( .A0(N132), .A1(N548), .B0(OFFSET[8]), .B1(N140), .Y(C2_Z_10) );
  AND2X2TF U151 ( .A(N345), .B(N223), .Y(N941) );
  AND2X2TF U152 ( .A(N354), .B(DP_OP_333_124_4748_N57), .Y(N747) );
  INVX1TF U153 ( .A(N345), .Y(N955) );
  OR2X2TF U154 ( .A(N169), .B(N246), .Y(N259) );
  OR2X2TF U155 ( .A(N351), .B(N600), .Y(N813) );
  AND2X2TF U156 ( .A(N123), .B(N246), .Y(N261) );
  NAND2XLTF U157 ( .A(N223), .B(N946), .Y(N534) );
  AND2X2TF U158 ( .A(N224), .B(ALU_START), .Y(N971) );
  CLKAND2X2TF U159 ( .A(ZTEMP[9]), .B(N142), .Y(POUT[9]) );
  CLKAND2X2TF U160 ( .A(ZTEMP[7]), .B(N142), .Y(POUT[7]) );
  CLKAND2X2TF U161 ( .A(ZTEMP[8]), .B(N142), .Y(POUT[8]) );
  AOI22X1TF U162 ( .A0(N73), .A1(DIVISION_HEAD[3]), .B0(XTEMP[12]), .B1(N61), 
        .Y(N349) );
  CLKAND2X2TF U163 ( .A(ZTEMP[10]), .B(N142), .Y(POUT[10]) );
  CLKAND2X2TF U164 ( .A(ZTEMP[12]), .B(N142), .Y(POUT[12]) );
  CLKINVX2TF U165 ( .A(N500), .Y(N82) );
  CLKAND2X2TF U166 ( .A(ZTEMP[11]), .B(N142), .Y(POUT[11]) );
  CLKAND2X2TF U167 ( .A(ZTEMP[1]), .B(N195), .Y(POUT[1]) );
  INVX2TF U168 ( .A(N200), .Y(N105) );
  CLKAND2X2TF U169 ( .A(ZTEMP[0]), .B(N195), .Y(POUT[0]) );
  CLKAND2X2TF U170 ( .A(ZTEMP[2]), .B(N195), .Y(POUT[2]) );
  AND2X1TF U171 ( .A(\INDEX[2] ), .B(N625), .Y(N314) );
  CLKAND2X2TF U172 ( .A(ZTEMP[5]), .B(N195), .Y(POUT[5]) );
  INVX2TF U173 ( .A(N73), .Y(N117) );
  CLKAND2X2TF U174 ( .A(ZTEMP[3]), .B(N195), .Y(POUT[3]) );
  INVX2TF U175 ( .A(N198), .Y(N89) );
  CLKAND2X2TF U176 ( .A(ZTEMP[4]), .B(N195), .Y(POUT[4]) );
  CLKAND2X2TF U177 ( .A(ZTEMP[6]), .B(N195), .Y(POUT[6]) );
  NAND2XLTF U178 ( .A(DIVISION_HEAD[4]), .B(N263), .Y(N226) );
  INVX2TF U179 ( .A(X_IN[5]), .Y(N200) );
  INVX2TF U180 ( .A(X_IN[11]), .Y(N201) );
  INVX2TF U181 ( .A(X_IN[3]), .Y(N199) );
  INVX2TF U182 ( .A(Y_IN[7]), .Y(N198) );
  INVX2TF U183 ( .A(ALU_TYPE[1]), .Y(N202) );
  INVX2TF U184 ( .A(N244), .Y(N83) );
  INVX2TF U185 ( .A(N244), .Y(N84) );
  INVX2TF U186 ( .A(N245), .Y(N85) );
  INVX2TF U187 ( .A(N245), .Y(N86) );
  INVX2TF U188 ( .A(N1019), .Y(N87) );
  INVX2TF U189 ( .A(N1019), .Y(N88) );
  INVX2TF U190 ( .A(N199), .Y(N93) );
  INVX2TF U191 ( .A(N199), .Y(N94) );
  INVX2TF U192 ( .A(N501), .Y(N95) );
  INVX2TF U193 ( .A(N501), .Y(N96) );
  INVX2TF U194 ( .A(N736), .Y(N98) );
  INVX2TF U195 ( .A(N747), .Y(N100) );
  INVX2TF U196 ( .A(N394), .Y(N101) );
  INVX2TF U197 ( .A(N394), .Y(N102) );
  INVX2TF U198 ( .A(N263), .Y(N103) );
  INVX2TF U199 ( .A(N263), .Y(N104) );
  INVX2TF U200 ( .A(N200), .Y(N106) );
  INVX2TF U201 ( .A(N1012), .Y(N107) );
  INVX2TF U202 ( .A(N1012), .Y(N108) );
  INVX2TF U203 ( .A(N259), .Y(N110) );
  INVX2TF U204 ( .A(N261), .Y(N111) );
  INVX2TF U205 ( .A(N261), .Y(N112) );
  INVX2TF U206 ( .A(N221), .Y(N113) );
  INVX2TF U207 ( .A(N221), .Y(N114) );
  INVX2TF U208 ( .A(N937), .Y(N115) );
  INVX2TF U209 ( .A(N937), .Y(N116) );
  INVX2TF U210 ( .A(N941), .Y(N119) );
  INVX2TF U211 ( .A(N813), .Y(N125) );
  INVX2TF U212 ( .A(N509), .Y(N126) );
  INVX2TF U213 ( .A(N509), .Y(N127) );
  INVX2TF U214 ( .A(N118), .Y(N130) );
  INVX2TF U215 ( .A(N97), .Y(N131) );
  INVX2TF U216 ( .A(N971), .Y(N132) );
  INVX2TF U217 ( .A(N971), .Y(N133) );
  AOI222X4TF U218 ( .A0(N487), .A1(N161), .B0(N487), .B1(N502), .C0(N161), 
        .C1(N502), .Y(N497) );
  NOR2X2TF U219 ( .A(N342), .B(N956), .Y(N354) );
  NOR3X2TF U220 ( .A(N118), .B(N605), .C(N632), .Y(N618) );
  INVX2TF U221 ( .A(N505), .Y(N134) );
  INVX2TF U222 ( .A(N505), .Y(N135) );
  INVX2TF U223 ( .A(N801), .Y(N136) );
  INVX2TF U224 ( .A(N801), .Y(N137) );
  NAND2X2TF U225 ( .A(N123), .B(N763), .Y(N454) );
  AOI21X2TF U226 ( .A0(N941), .A1(N921), .B0(N222), .Y(N935) );
  INVX2TF U227 ( .A(N201), .Y(N138) );
  INVX2TF U228 ( .A(N201), .Y(N139) );
  AOI211XLTF U229 ( .A0(N832), .A1(N831), .B0(OPER_A[2]), .C0(N916), .Y(N833)
         );
  OAI32XLTF U230 ( .A0(OPER_A[8]), .A1(N898), .A2(N916), .B0(N897), .B1(N896), 
        .Y(N899) );
  OAI32XLTF U231 ( .A0(OPER_A[10]), .A1(N917), .A2(N916), .B0(N915), .B1(N914), 
        .Y(N918) );
  OAI32XLTF U232 ( .A0(OPER_A[6]), .A1(N882), .A2(N916), .B0(N881), .B1(N880), 
        .Y(N883) );
  INVXLTF U233 ( .A(N916), .Y(N913) );
  INVXLTF U234 ( .A(X_IN[2]), .Y(N772) );
  INVX2TF U235 ( .A(DP_OP_333_124_4748_N57), .Y(N140) );
  INVX2TF U236 ( .A(N969), .Y(N141) );
  AOI2BB1X2TF U237 ( .A0N(N963), .A1N(N962), .B0(N961), .Y(N1011) );
  CLKBUFX2TF U238 ( .A(N195), .Y(N142) );
  CLKBUFX2TF U239 ( .A(N262), .Y(N195) );
  NOR3XLTF U240 ( .A(N73), .B(N910), .C(N972), .Y(N821) );
  NAND2X2TF U241 ( .A(N970), .B(N929), .Y(N910) );
  AOI21XLTF U242 ( .A0(N824), .A1(N823), .B0(N822), .Y(N835) );
  INVXLTF U243 ( .A(N822), .Y(N379) );
  NOR3BX4TF U244 ( .AN(N384), .B(N381), .C(N131), .Y(N513) );
  AOI222X4TF U245 ( .A0(XTEMP[9]), .A1(X_IN[9]), .B0(XTEMP[9]), .B1(N478), 
        .C0(X_IN[9]), .C1(N478), .Y(N487) );
  AOI222X4TF U246 ( .A0(N178), .A1(N488), .B0(N178), .B1(N464), .C0(N488), 
        .C1(N464), .Y(N478) );
  OAI31XLTF U247 ( .A0(OPER_A[1]), .A1(N916), .A2(OPER_A[0]), .B0(N837), .Y(
        N838) );
  OAI21X2TF U248 ( .A0(N514), .A1(N111), .B0(N248), .Y(OPER_A[1]) );
  INVX2TF U249 ( .A(N123), .Y(N143) );
  NAND2X2TF U250 ( .A(N763), .B(N143), .Y(N559) );
  AOI22XLTF U251 ( .A0(X_IN[1]), .A1(N807), .B0(X_IN[0]), .B1(N136), .Y(N754)
         );
  AOI22XLTF U252 ( .A0(X_IN[4]), .A1(N101), .B0(X_IN[6]), .B1(N807), .Y(N552)
         );
  AOI22XLTF U253 ( .A0(X_IN[12]), .A1(N807), .B0(N139), .B1(N136), .Y(N436) );
  AOI22XLTF U254 ( .A0(X_IN[2]), .A1(N101), .B0(X_IN[4]), .B1(N807), .Y(N792)
         );
  AOI22XLTF U255 ( .A0(DIVISION_HEAD[5]), .A1(N95), .B0(X_IN[7]), .B1(N807), 
        .Y(N387) );
  AOI22XLTF U256 ( .A0(X_IN[10]), .A1(N136), .B0(N139), .B1(N807), .Y(N427) );
  AOI22XLTF U257 ( .A0(X_IN[2]), .A1(N136), .B0(N94), .B1(N807), .Y(N786) );
  AOI22XLTF U258 ( .A0(N94), .A1(N101), .B0(N106), .B1(N807), .Y(N808) );
  NOR4X2TF U259 ( .A(N648), .B(N943), .C(N370), .D(N369), .Y(N642) );
  NOR2X2TF U260 ( .A(N342), .B(N604), .Y(N566) );
  NOR2BX2TF U261 ( .AN(N544), .B(N382), .Y(N629) );
  NOR2X2TF U262 ( .A(N351), .B(N132), .Y(N382) );
  INVX2TF U263 ( .A(N144), .Y(N145) );
  INVX2TF U264 ( .A(N144), .Y(N146) );
  AOI22X2TF U265 ( .A0(N349), .A1(N347), .B0(N940), .B1(N350), .Y(N922) );
  NOR3X4TF U266 ( .A(N202), .B(ALU_TYPE[0]), .C(ALU_TYPE[2]), .Y(N224) );
  XNOR2X1TF U267 ( .A(OPER_A[12]), .B(ADD_X_132_1_N2), .Y(N147) );
  XNOR2X2TF U268 ( .A(N147), .B(OPER_B[12]), .Y(SUM_AB[12]) );
  ADDHX1TF U269 ( .A(OPER_B[0]), .B(OPER_A[0]), .CO(ADD_X_132_1_N13), .S(
        SUM_AB[0]) );
  INVX2TF U270 ( .A(OPER_A[0]), .Y(N831) );
  AOI222XLTF U271 ( .A0(DIVISION_HEAD[1]), .A1(DIVISION_HEAD[0]), .B0(
        DIVISION_HEAD[1]), .B1(N318), .C0(DIVISION_HEAD[0]), .C1(N317), .Y(
        N320) );
  AOI32X1TF U272 ( .A0(N941), .A1(N61), .A2(N564), .B0(N618), .B1(N73), .Y(
        N545) );
  AOI22X1TF U273 ( .A0(N73), .A1(N167), .B0(POST_WORK), .B1(N117), .Y(N246) );
  OAI31X1TF U274 ( .A0(N133), .A1(N949), .A2(N948), .B0(N947), .Y(N950) );
  NAND2X1TF U275 ( .A(N317), .B(N727), .Y(N319) );
  INVX2TF U276 ( .A(N929), .Y(N222) );
  OAI21X1TF U277 ( .A0(N948), .A1(N610), .B0(N647), .Y(N961) );
  NAND2X1TF U278 ( .A(N477), .B(N476), .Y(N486) );
  NOR2X1TF U279 ( .A(SUM_AB[8]), .B(N462), .Y(N477) );
  OA22X1TF U280 ( .A0(N769), .A1(N558), .B0(N764), .B1(N765), .Y(N309) );
  NOR2X2TF U281 ( .A(N222), .B(N118), .Y(N904) );
  OR2X2TF U282 ( .A(N961), .B(N203), .Y(N929) );
  OAI21X1TF U283 ( .A0(DIVISION_HEAD[12]), .A1(N549), .B0(N341), .Y(N948) );
  AOI2BB1X1TF U284 ( .A0N(DIVISION_HEAD[6]), .A1N(N330), .B0(Y_IN[6]), .Y(N328) );
  AOI21X1TF U285 ( .A0(N197), .A1(N514), .B0(N327), .Y(N330) );
  AOI2BB1X1TF U286 ( .A0N(DIVISION_HEAD[4]), .A1N(N326), .B0(Y_IN[4]), .Y(N324) );
  NOR2X1TF U287 ( .A(SUM_AB[10]), .B(N486), .Y(N499) );
  NOR2X1TF U288 ( .A(\INDEX[2] ), .B(N621), .Y(N312) );
  NAND2X1TF U289 ( .A(N129), .B(N128), .Y(N621) );
  NAND2X1TF U290 ( .A(N912), .B(N904), .Y(N932) );
  NAND2X1TF U291 ( .A(N565), .B(N350), .Y(N916) );
  AOI2BB1X1TF U292 ( .A0N(N608), .A1N(N346), .B0(N962), .Y(N203) );
  NAND2X1TF U293 ( .A(N566), .B(N382), .Y(N610) );
  AOI211X1TF U294 ( .A0(Y_IN[11]), .A1(N305), .B0(Y_IN[12]), .C0(N287), .Y(
        N767) );
  NOR2X1TF U295 ( .A(PRE_WORK), .B(N343), .Y(N345) );
  NOR2X1TF U296 ( .A(N124), .B(N628), .Y(N343) );
  NAND2X1TF U297 ( .A(N122), .B(N152), .Y(N605) );
  NAND2X1TF U298 ( .A(N180), .B(N368), .Y(N351) );
  NAND2X1TF U299 ( .A(N151), .B(N153), .Y(N342) );
  NAND2X1TF U300 ( .A(N454), .B(N460), .Y(N471) );
  NAND2X2TF U301 ( .A(N547), .B(N384), .Y(N460) );
  NAND2X1TF U302 ( .A(N121), .B(N170), .Y(N604) );
  CLKBUFX2TF U303 ( .A(N782), .Y(N196) );
  NAND2X1TF U304 ( .A(N121), .B(N122), .Y(N956) );
  NAND3X1TF U305 ( .A(N962), .B(N132), .C(N600), .Y(N647) );
  CLKBUFX2TF U306 ( .A(Y_IN[5]), .Y(N197) );
  AND2X2TF U307 ( .A(ALU_START), .B(N142), .Y(N223) );
  NAND2X1TF U308 ( .A(N124), .B(N312), .Y(N368) );
  NOR3X1TF U309 ( .A(N606), .B(N605), .C(N777), .Y(N607) );
  OR3X1TF U310 ( .A(N888), .B(N887), .C(N217), .Y(N676) );
  OAI2BB2XLTF U311 ( .B0(N889), .B1(N972), .A0N(C152_DATA4_6), .A1N(N114), .Y(
        N217) );
  OAI2BB2XLTF U312 ( .B0(N886), .B1(N924), .A0N(N222), .A1N(OPER_B[6]), .Y(
        N887) );
  AOI32X1TF U313 ( .A0(N970), .A1(N969), .A2(N968), .B0(N130), .B1(N969), .Y(
        N1019) );
  INVX2TF U314 ( .A(N460), .Y(N475) );
  NAND2X1TF U315 ( .A(N647), .B(N99), .Y(N944) );
  NAND2X1TF U316 ( .A(N566), .B(DP_OP_333_124_4748_N57), .Y(N393) );
  NAND2X1TF U317 ( .A(SIGN_Y), .B(N965), .Y(N972) );
  NAND2X1TF U318 ( .A(N904), .B(N877), .Y(N894) );
  INVX2TF U319 ( .A(DP_OP_333_124_4748_N57), .Y(N207) );
  AOI21X1TF U320 ( .A0(N949), .A1(N967), .B0(N366), .Y(N970) );
  NOR2BX2TF U321 ( .AN(N547), .B(N557), .Y(N814) );
  NAND2X1TF U322 ( .A(N151), .B(STEP[3]), .Y(N632) );
  NOR2X1TF U323 ( .A(N180), .B(N600), .Y(N356) );
  INVX2TF U324 ( .A(N223), .Y(N962) );
  NAND2X1TF U325 ( .A(N960), .B(DP_OP_333_124_4748_N57), .Y(N651) );
  AND2X2TF U326 ( .A(N223), .B(PRE_WORK), .Y(DP_OP_333_124_4748_N57) );
  INVX2TF U327 ( .A(N367), .Y(N763) );
  NAND2X1TF U328 ( .A(N382), .B(N960), .Y(N367) );
  NOR2X2TF U329 ( .A(N342), .B(N605), .Y(N960) );
  AO22X1TF U330 ( .A0(N375), .A1(XTEMP[12]), .B0(N363), .B1(N965), .Y(N722) );
  AOI211X1TF U331 ( .A0(N223), .A1(N608), .B0(N945), .C0(N607), .Y(N611) );
  AOI32X1TF U332 ( .A0(N967), .A1(N364), .A2(N958), .B0(N973), .B1(N364), .Y(
        N365) );
  NAND2X1TF U333 ( .A(N643), .B(N125), .Y(N615) );
  NAND2X1TF U334 ( .A(N946), .B(DP_OP_333_124_4748_N57), .Y(N635) );
  NAND2X1TF U335 ( .A(N114), .B(C152_DATA4_8), .Y(N218) );
  AOI32X1TF U336 ( .A0(N126), .A1(DIVISION_HEAD[4]), .A2(N750), .B0(N471), 
        .B1(DIVISION_HEAD[4]), .Y(N391) );
  OAI22X1TF U337 ( .A0(N529), .A1(N98), .B0(N488), .B1(N100), .Y(N489) );
  OAI22X1TF U338 ( .A0(N514), .A1(N97), .B0(N157), .B1(N454), .Y(N405) );
  OAI2BB2XLTF U339 ( .B0(N61), .B1(N972), .A0N(N972), .A1N(N61), .Y(N974) );
  OAI22X1TF U340 ( .A0(N161), .A1(N97), .B0(N500), .B1(N99), .Y(N504) );
  NAND2X1TF U341 ( .A(N132), .B(N140), .Y(N208) );
  NOR2X1TF U342 ( .A(N605), .B(N954), .Y(N565) );
  NAND2X1TF U343 ( .A(STEP[2]), .B(N153), .Y(N954) );
  INVX2TF U344 ( .A(N120), .Y(N777) );
  NOR2X2TF U345 ( .A(N763), .B(N196), .Y(N761) );
  NAND2X1TF U346 ( .A(N354), .B(N120), .Y(N544) );
  NOR2X1TF U347 ( .A(N956), .B(N632), .Y(N564) );
  OAI21X2TF U348 ( .A0(N158), .A1(N111), .B0(N247), .Y(OPER_A[0]) );
  OAI32X1TF U349 ( .A0(N650), .A1(N182), .A2(N944), .B0(N649), .B1(N651), .Y(
        N694) );
  OAI21X1TF U350 ( .A0(N180), .A1(N648), .B0(N647), .Y(N695) );
  AOI22X1TF U351 ( .A0(N543), .A1(N73), .B0(N542), .B1(N541), .Y(N707) );
  INVX2TF U352 ( .A(N543), .Y(N541) );
  OAI31X1TF U353 ( .A0(N540), .A1(N539), .A2(N538), .B0(N537), .Y(N542) );
  AOI211X1TF U354 ( .A0(N536), .A1(XTEMP[12]), .B0(N535), .C0(N534), .Y(N537)
         );
  OAI31X1TF U355 ( .A0(DIVISION_HEAD[1]), .A1(N533), .A2(N161), .B0(N532), .Y(
        N536) );
  AOI22X1TF U356 ( .A0(N531), .A1(N530), .B0(XTEMP[11]), .B1(N168), .Y(N532)
         );
  OAI22X1TF U357 ( .A0(DIVISION_HEAD[0]), .A1(N529), .B0(DIVISION_REMA[8]), 
        .B1(N178), .Y(N530) );
  INVX2TF U358 ( .A(N539), .Y(N531) );
  NOR2X1TF U359 ( .A(XTEMP[11]), .B(N168), .Y(N533) );
  OAI22X1TF U360 ( .A0(DIVISION_HEAD[12]), .A1(N149), .B0(XTEMP[12]), .B1(N649), .Y(N538) );
  OAI21X1TF U361 ( .A0(XTEMP[11]), .A1(N168), .B0(N528), .Y(N539) );
  AOI22X1TF U362 ( .A0(DIVISION_HEAD[0]), .A1(N529), .B0(DIVISION_HEAD[1]), 
        .B1(N161), .Y(N528) );
  AOI21X1TF U363 ( .A0(DIVISION_HEAD[11]), .A1(N173), .B0(N527), .Y(N540) );
  AOI211X1TF U364 ( .A0(DIVISION_REMA[6]), .A1(N160), .B0(N526), .C0(N525), 
        .Y(N527) );
  NOR2X1TF U365 ( .A(DIVISION_HEAD[11]), .B(N173), .Y(N525) );
  AOI21X1TF U366 ( .A0(DIVISION_HEAD[9]), .A1(N172), .B0(N523), .Y(N524) );
  AOI211X1TF U367 ( .A0(DIVISION_REMA[4]), .A1(N155), .B0(N522), .C0(N521), 
        .Y(N523) );
  NOR2X1TF U368 ( .A(DIVISION_HEAD[9]), .B(N172), .Y(N521) );
  AOI21X1TF U369 ( .A0(DIVISION_HEAD[7]), .A1(N171), .B0(N519), .Y(N520) );
  AOI211X1TF U370 ( .A0(N518), .A1(DIVISION_REMA[2]), .B0(N517), .C0(N516), 
        .Y(N519) );
  NOR2X1TF U371 ( .A(DIVISION_HEAD[7]), .B(N171), .Y(N517) );
  OAI21X1TF U372 ( .A0(DIVISION_HEAD[5]), .A1(N184), .B0(N515), .Y(N518) );
  OAI211X1TF U373 ( .A0(DIVISION_REMA[1]), .A1(N514), .B0(DIVISION_REMA[0]), 
        .C0(N158), .Y(N515) );
  OAI21X1TF U374 ( .A0(N123), .A1(N952), .B0(N951), .Y(N670) );
  OAI21X1TF U375 ( .A0(N950), .A1(N970), .B0(N952), .Y(N951) );
  OR4X2TF U376 ( .A(N945), .B(N944), .C(N943), .D(N942), .Y(N952) );
  OAI22X1TF U377 ( .A0(N119), .A1(N940), .B0(N939), .B1(N973), .Y(N942) );
  OAI21X1TF U378 ( .A0(N597), .A1(N586), .B0(N585), .Y(N702) );
  AOI31X1TF U379 ( .A0(N584), .A1(N589), .A2(N591), .B0(N583), .Y(N586) );
  OAI22X1TF U380 ( .A0(N128), .A1(N582), .B0(N593), .B1(N589), .Y(N583) );
  OAI21X1TF U381 ( .A0(N128), .A1(N620), .B0(N619), .Y(N699) );
  AOI31X1TF U382 ( .A0(N618), .A1(N621), .A2(N617), .B0(N616), .Y(N619) );
  OAI32X1TF U383 ( .A0(N629), .A1(N630), .A2(N621), .B0(N617), .B1(N629), .Y(
        N616) );
  AOI22X1TF U384 ( .A0(N597), .A1(N92), .B0(N581), .B1(N580), .Y(N703) );
  AOI211X1TF U385 ( .A0(N595), .A1(N163), .B0(N579), .C0(N791), .Y(N581) );
  AOI21X1TF U386 ( .A0(N578), .A1(N777), .B0(N185), .Y(N579) );
  OAI31X1TF U387 ( .A0(N630), .A1(N629), .A2(N628), .B0(N627), .Y(N698) );
  AOI22X1TF U388 ( .A0(\INDEX[2] ), .A1(N626), .B0(N625), .B1(N624), .Y(N627)
         );
  OAI21X1TF U389 ( .A0(N623), .A1(N629), .B0(N622), .Y(N626) );
  OAI211X1TF U390 ( .A0(N119), .A1(N372), .B0(N645), .C0(N371), .Y(N721) );
  AOI22X1TF U391 ( .A0(STEP[3]), .A1(N642), .B0(N377), .B1(N574), .Y(N371) );
  OAI211X1TF U392 ( .A0(N183), .A1(N615), .B0(N631), .C0(N614), .Y(N700) );
  AOI21X1TF U393 ( .A0(N642), .A1(N152), .B0(N613), .Y(N614) );
  NOR3X1TF U394 ( .A(STEP[3]), .B(N119), .C(N604), .Y(N945) );
  AOI211X1TF U395 ( .A0(N824), .A1(N377), .B0(N375), .C0(N374), .Y(N612) );
  AOI21X1TF U396 ( .A0(N383), .A1(N373), .B0(N777), .Y(N374) );
  NOR2X1TF U397 ( .A(N118), .B(N823), .Y(N377) );
  OAI22X1TF U398 ( .A0(N90), .A1(N598), .B0(N597), .B1(N596), .Y(N701) );
  AOI21X1TF U399 ( .A0(\INDEX[2] ), .A1(N595), .B0(N594), .Y(N596) );
  OAI22X1TF U400 ( .A0(N593), .A1(N592), .B0(N591), .B1(N590), .Y(N594) );
  INVX2TF U401 ( .A(N588), .Y(N593) );
  AOI21X1TF U402 ( .A0(N589), .A1(N588), .B0(N587), .Y(N598) );
  OAI211X1TF U403 ( .A0(N646), .A1(N151), .B0(N645), .C0(N644), .Y(N696) );
  NOR2X1TF U404 ( .A(N650), .B(N365), .Y(N645) );
  INVX2TF U405 ( .A(N651), .Y(N650) );
  OAI22X1TF U406 ( .A0(N170), .A1(N954), .B0(N823), .B1(N967), .Y(N638) );
  AOI211X1TF U407 ( .A0(N642), .A1(N170), .B0(N637), .C0(N636), .Y(N641) );
  AOI21X1TF U408 ( .A0(N81), .A1(N603), .B0(N602), .Y(N631) );
  OAI21X1TF U409 ( .A0(N601), .A1(N600), .B0(N599), .Y(N602) );
  OAI22X1TF U410 ( .A0(N597), .A1(N577), .B0(N576), .B1(N194), .Y(N704) );
  AOI21X1TF U411 ( .A0(N592), .A1(N588), .B0(N587), .Y(N576) );
  OAI21X1TF U412 ( .A0(N90), .A1(N591), .B0(N584), .Y(N590) );
  INVX2TF U413 ( .A(N615), .Y(N584) );
  INVX2TF U414 ( .A(N597), .Y(N580) );
  OAI31X1TF U415 ( .A0(N606), .A1(N605), .A2(N777), .B0(N578), .Y(N588) );
  OAI32X1TF U416 ( .A0(N575), .A1(N824), .A2(N574), .B0(N130), .B1(N575), .Y(
        N578) );
  INVX2TF U417 ( .A(N573), .Y(N575) );
  AOI21X1TF U418 ( .A0(N595), .A1(N191), .B0(N572), .Y(N577) );
  AOI32X1TF U419 ( .A0(N566), .A1(N125), .A2(N183), .B0(N960), .B1(N120), .Y(
        N568) );
  AOI31X1TF U420 ( .A0(N130), .A1(N824), .A2(N823), .B0(N944), .Y(N569) );
  INVX2TF U421 ( .A(N582), .Y(N595) );
  AOI32X1TF U422 ( .A0(N314), .A1(N124), .A2(N618), .B0(N191), .B1(N313), .Y(
        N316) );
  NOR2X1TF U423 ( .A(N630), .B(N624), .Y(N622) );
  AOI21X1TF U424 ( .A0(\INDEX[2] ), .A1(N625), .B0(N378), .Y(N624) );
  INVX2TF U425 ( .A(N620), .Y(N630) );
  INVX2TF U426 ( .A(N617), .Y(N625) );
  OAI21X1TF U427 ( .A0(N129), .A1(N620), .B0(N311), .Y(N726) );
  OAI21X1TF U428 ( .A0(N310), .A1(N381), .B0(N620), .Y(N311) );
  AOI32X1TF U429 ( .A0(N629), .A1(N635), .A2(N378), .B0(N163), .B1(N635), .Y(
        N310) );
  INVX2TF U430 ( .A(N265), .Y(N634) );
  AOI31X1TF U431 ( .A0(N956), .A1(N373), .A2(N383), .B0(N777), .Y(N265) );
  OAI21X1TF U432 ( .A0(N354), .A1(N264), .B0(N941), .Y(N364) );
  AOI22X1TF U433 ( .A0(N903), .A1(N904), .B0(N222), .B1(OPER_B[8]), .Y(N219)
         );
  OAI21X1TF U434 ( .A0(N902), .A1(N165), .B0(N901), .Y(N903) );
  AOI211X1TF U435 ( .A0(N920), .A1(OPER_B[9]), .B0(N900), .C0(N899), .Y(N901)
         );
  AOI21X1TF U436 ( .A0(N913), .A1(N898), .B0(N912), .Y(N896) );
  NOR3X1TF U437 ( .A(N911), .B(OPER_B[8]), .C(N895), .Y(N900) );
  AOI21X1TF U438 ( .A0(N895), .A1(N922), .B0(N921), .Y(N902) );
  INVX2TF U439 ( .A(N888), .Y(N214) );
  AOI31X1TF U440 ( .A0(N842), .A1(N841), .A2(N840), .B0(N924), .Y(N844) );
  AOI32X1TF U441 ( .A0(N839), .A1(OPER_B[2]), .A2(N922), .B0(N921), .B1(
        OPER_B[2]), .Y(N840) );
  AOI22X1TF U442 ( .A0(N920), .A1(OPER_B[3]), .B0(OPER_A[2]), .B1(N838), .Y(
        N841) );
  AOI31X1TF U443 ( .A0(N922), .A1(N162), .A2(N834), .B0(N833), .Y(N842) );
  OAI211X1TF U444 ( .A0(N1010), .A1(N997), .B0(N996), .C0(N995), .Y(N662) );
  AOI22X1TF U445 ( .A0(DIVISION_HEAD[7]), .A1(N107), .B0(ZTEMP[7]), .B1(N141), 
        .Y(N996) );
  OAI211X1TF U446 ( .A0(N1010), .A1(N1003), .B0(N1002), .C0(N1001), .Y(N660)
         );
  AOI22X1TF U447 ( .A0(DIVISION_HEAD[9]), .A1(N107), .B0(ZTEMP[9]), .B1(N1011), 
        .Y(N1002) );
  OAI211X1TF U448 ( .A0(N1010), .A1(N991), .B0(N990), .C0(N989), .Y(N664) );
  AOI22X1TF U449 ( .A0(DIVISION_HEAD[5]), .A1(N107), .B0(ZTEMP[5]), .B1(N141), 
        .Y(N990) );
  OAI211X1TF U450 ( .A0(N1010), .A1(N985), .B0(N984), .C0(N983), .Y(N666) );
  AOI22X1TF U451 ( .A0(DIVISION_HEAD[3]), .A1(N107), .B0(ZTEMP[3]), .B1(N1011), 
        .Y(N984) );
  AOI211X1TF U452 ( .A0(N222), .A1(OPER_B[10]), .B0(N927), .C0(N928), .Y(N220)
         );
  AOI21X1TF U453 ( .A0(N975), .A1(N972), .B0(N910), .Y(N928) );
  AOI21X1TF U454 ( .A0(N926), .A1(N925), .B0(N924), .Y(N927) );
  AOI32X1TF U455 ( .A0(N923), .A1(OPER_B[10]), .A2(N922), .B0(N921), .B1(
        OPER_B[10]), .Y(N925) );
  AOI211X1TF U456 ( .A0(N920), .A1(OPER_B[11]), .B0(N919), .C0(N918), .Y(N926)
         );
  AOI21X1TF U457 ( .A0(N913), .A1(N917), .B0(N912), .Y(N914) );
  NOR3X1TF U458 ( .A(N911), .B(OPER_B[10]), .C(N923), .Y(N919) );
  AOI22X1TF U459 ( .A0(SUM_AB[2]), .A1(N87), .B0(N980), .B1(N1015), .Y(N981)
         );
  AOI22X1TF U460 ( .A0(DIVISION_HEAD[2]), .A1(N108), .B0(ZTEMP[2]), .B1(N141), 
        .Y(N982) );
  AOI22X1TF U461 ( .A0(SUM_AB[1]), .A1(N87), .B0(N977), .B1(N1015), .Y(N978)
         );
  AOI22X1TF U462 ( .A0(DIVISION_HEAD[1]), .A1(N108), .B0(ZTEMP[1]), .B1(N141), 
        .Y(N979) );
  AOI22X1TF U463 ( .A0(SUM_AB[6]), .A1(N87), .B0(N992), .B1(N1015), .Y(N993)
         );
  AOI22X1TF U464 ( .A0(DIVISION_HEAD[6]), .A1(N108), .B0(ZTEMP[6]), .B1(N141), 
        .Y(N994) );
  AOI22X1TF U465 ( .A0(SUM_AB[4]), .A1(N87), .B0(N986), .B1(N1015), .Y(N987)
         );
  AOI22X1TF U466 ( .A0(DIVISION_HEAD[4]), .A1(N108), .B0(ZTEMP[4]), .B1(N141), 
        .Y(N988) );
  AOI22X1TF U467 ( .A0(SUM_AB[8]), .A1(N87), .B0(N998), .B1(N1015), .Y(N999)
         );
  AOI22X1TF U468 ( .A0(DIVISION_HEAD[8]), .A1(N108), .B0(ZTEMP[8]), .B1(N141), 
        .Y(N1000) );
  AOI211X1TF U469 ( .A0(OPER_B[6]), .A1(N885), .B0(N884), .C0(N883), .Y(N886)
         );
  AOI21X1TF U470 ( .A0(N913), .A1(N882), .B0(N912), .Y(N880) );
  OAI31X1TF U471 ( .A0(N911), .A1(OPER_B[6]), .A2(N879), .B0(N878), .Y(N884)
         );
  AOI21X1TF U472 ( .A0(OPER_B[7]), .A1(N877), .B0(N876), .Y(N878) );
  OAI21X1TF U473 ( .A0(N911), .A1(N875), .B0(N874), .Y(N885) );
  OAI22X1TF U474 ( .A0(N475), .A1(N474), .B0(N473), .B1(N178), .Y(N711) );
  AOI211X1TF U475 ( .A0(N998), .A1(N493), .B0(N470), .C0(N469), .Y(N474) );
  OAI211X1TF U476 ( .A0(N468), .A1(N609), .B0(N467), .C0(N466), .Y(N469) );
  AOI22X1TF U477 ( .A0(XTEMP[9]), .A1(N96), .B0(N800), .B1(SUM_AB[12]), .Y(
        N466) );
  NOR2X1TF U478 ( .A(DIVISION_HEAD[12]), .B(N472), .Y(N465) );
  AOI22X1TF U479 ( .A0(X_IN[8]), .A1(N464), .B0(INTADD_0_N1), .B1(N488), .Y(
        N472) );
  OAI22X1TF U480 ( .A0(N154), .A1(N98), .B0(N463), .B1(N100), .Y(N470) );
  AOI22X1TF U481 ( .A0(SUM_AB[10]), .A1(N88), .B0(N1004), .B1(N1015), .Y(N1005) );
  AOI22X1TF U482 ( .A0(DIVISION_HEAD[10]), .A1(N108), .B0(ZTEMP[10]), .B1(N141), .Y(N1006) );
  OAI21X1TF U483 ( .A0(N450), .A1(N449), .B0(N460), .Y(N451) );
  AOI22X1TF U484 ( .A0(DIVISION_HEAD[11]), .A1(N96), .B0(X_IN[12]), .B1(N137), 
        .Y(N445) );
  AOI22X1TF U485 ( .A0(N106), .A1(N444), .B0(N139), .B1(N102), .Y(N446) );
  AOI22X1TF U486 ( .A0(SUM_AB[6]), .A1(N134), .B0(N493), .B1(N992), .Y(N447)
         );
  OAI22X1TF U487 ( .A0(N156), .A1(N98), .B0(N442), .B1(N100), .Y(N450) );
  AOI32X1TF U488 ( .A0(N431), .A1(N460), .A2(N430), .B0(N475), .B1(N155), .Y(
        N715) );
  AOI211X1TF U489 ( .A0(N493), .A1(N986), .B0(N429), .C0(N428), .Y(N430) );
  AOI22X1TF U490 ( .A0(DIVISION_HEAD[9]), .A1(N95), .B0(N82), .B1(N102), .Y(
        N426) );
  OAI22X1TF U491 ( .A0(N423), .A1(N98), .B0(N155), .B1(N454), .Y(N429) );
  AOI32X1TF U492 ( .A0(N392), .A1(N391), .A2(N390), .B0(N475), .B1(N391), .Y(
        N719) );
  OAI211X1TF U493 ( .A0(N388), .A1(N559), .B0(N387), .C0(N386), .Y(N389) );
  AOI22X1TF U494 ( .A0(X_IN[6]), .A1(N137), .B0(N106), .B1(N102), .Y(N386) );
  AOI22X1TF U495 ( .A0(DIVISION_HEAD[3]), .A1(N736), .B0(SUM_AB[0]), .B1(N380), 
        .Y(N392) );
  AOI32X1TF U496 ( .A0(N401), .A1(N460), .A2(N400), .B0(N475), .B1(N514), .Y(
        N718) );
  AOI211X1TF U497 ( .A0(N493), .A1(N977), .B0(N399), .C0(N398), .Y(N400) );
  OAI211X1TF U498 ( .A0(N559), .A1(N432), .B0(N397), .C0(N396), .Y(N398) );
  AOI21X1TF U499 ( .A0(DIVISION_HEAD[4]), .A1(N736), .B0(N395), .Y(N396) );
  OAI22X1TF U500 ( .A0(N514), .A1(N454), .B0(N750), .B1(N609), .Y(N395) );
  AOI22X1TF U501 ( .A0(DIVISION_HEAD[6]), .A1(N96), .B0(X_IN[7]), .B1(N137), 
        .Y(N397) );
  OAI22X1TF U502 ( .A0(N463), .A1(N394), .B0(N488), .B1(N749), .Y(N399) );
  OAI22X1TF U503 ( .A0(N513), .A1(N496), .B0(N495), .B1(N161), .Y(N709) );
  AOI21X1TF U504 ( .A0(N493), .A1(N1004), .B0(N492), .Y(N496) );
  OAI211X1TF U505 ( .A0(N500), .A1(N609), .B0(N491), .C0(N490), .Y(N492) );
  AOI22X1TF U506 ( .A0(XTEMP[11]), .A1(N96), .B0(SUM_AB[10]), .B1(N134), .Y(
        N491) );
  AOI32X1TF U507 ( .A0(N411), .A1(N460), .A2(N410), .B0(N475), .B1(N157), .Y(
        N717) );
  AOI211X1TF U508 ( .A0(DIVISION_HEAD[7]), .A1(N96), .B0(N409), .C0(N408), .Y(
        N410) );
  OAI211X1TF U509 ( .A0(N100), .A1(N750), .B0(N407), .C0(N406), .Y(N408) );
  AOI21X1TF U510 ( .A0(N493), .A1(N980), .B0(N405), .Y(N406) );
  AOI22X1TF U511 ( .A0(X_IN[1]), .A1(N444), .B0(N800), .B1(SUM_AB[6]), .Y(N407) );
  OAI21X1TF U512 ( .A0(N500), .A1(N749), .B0(N402), .Y(N409) );
  AOI22X1TF U513 ( .A0(X_IN[8]), .A1(N137), .B0(X_IN[7]), .B1(N102), .Y(N402)
         );
  OAI211X1TF U514 ( .A0(N1010), .A1(N1009), .B0(N1008), .C0(N1007), .Y(N658)
         );
  AOI22X1TF U515 ( .A0(DIVISION_HEAD[11]), .A1(N108), .B0(ZTEMP[11]), .B1(N141), .Y(N1008) );
  INVX2TF U516 ( .A(N1015), .Y(N1010) );
  OAI211X1TF U517 ( .A0(N1019), .A1(N1018), .B0(N1017), .C0(N1016), .Y(N657)
         );
  AOI32X1TF U518 ( .A0(N1018), .A1(N1015), .A2(N1014), .B0(N1013), .B1(N1015), 
        .Y(N1016) );
  AOI211X4TF U519 ( .A0(N975), .A1(N974), .B0(N973), .C0(N1011), .Y(N1015) );
  INVX2TF U520 ( .A(N970), .Y(N973) );
  AOI22X1TF U521 ( .A0(DIVISION_HEAD[12]), .A1(N108), .B0(ZTEMP[12]), .B1(
        N1011), .Y(N1017) );
  OAI31X1TF U522 ( .A0(N967), .A1(N61), .A2(N972), .B0(N966), .Y(N968) );
  AOI31X1TF U523 ( .A0(N182), .A1(N61), .A2(N965), .B0(N964), .Y(N966) );
  INVX2TF U524 ( .A(N1011), .Y(N969) );
  AOI31X1TF U525 ( .A0(N960), .A1(N959), .A2(N958), .B0(N957), .Y(N963) );
  OAI31X1TF U526 ( .A0(N956), .A1(N955), .A2(N954), .B0(N953), .Y(N957) );
  INVX2TF U527 ( .A(N922), .Y(N911) );
  OAI22X1TF U528 ( .A0(N513), .A1(N512), .B0(N511), .B1(N159), .Y(N708) );
  OAI21X1TF U529 ( .A0(N507), .A1(N1009), .B0(N506), .Y(N508) );
  AOI211X1TF U530 ( .A0(SUM_AB[11]), .A1(N134), .B0(N504), .C0(N503), .Y(N506)
         );
  OAI22X1TF U531 ( .A0(N513), .A1(N485), .B0(N484), .B1(N529), .Y(N710) );
  AOI211X1TF U532 ( .A0(SUM_AB[9]), .A1(N135), .B0(N482), .C0(N481), .Y(N485)
         );
  OAI211X1TF U533 ( .A0(N1003), .A1(N507), .B0(N480), .C0(N479), .Y(N481) );
  OAI22X1TF U534 ( .A0(N178), .A1(N98), .B0(N488), .B1(N609), .Y(N482) );
  AOI32X1TF U535 ( .A0(N799), .A1(N816), .A2(N798), .B0(N814), .B1(N175), .Y(
        N684) );
  AOI21X1TF U536 ( .A0(N797), .A1(N1004), .B0(N796), .Y(N798) );
  AOI22X1TF U537 ( .A0(DIVISION_HEAD[0]), .A1(N131), .B0(DIVISION_HEAD[1]), 
        .B1(N806), .Y(N793) );
  AOI22X1TF U538 ( .A0(Y_IN[10]), .A1(N791), .B0(N94), .B1(N137), .Y(N794) );
  AOI21X1TF U539 ( .A0(SUM_AB[10]), .A1(N486), .B0(N499), .Y(N1004) );
  AOI22X1TF U540 ( .A0(N800), .A1(SUM_AB[1]), .B0(SUM_AB[10]), .B1(N146), .Y(
        N799) );
  OAI21X1TF U541 ( .A0(N761), .A1(N183), .B0(N563), .Y(N705) );
  OAI22X1TF U542 ( .A0(N562), .A1(N561), .B0(N763), .B1(N780), .Y(N563) );
  AOI22X1TF U543 ( .A0(Y_IN[0]), .A1(N791), .B0(DIVISION_REMA[1]), .B1(N120), 
        .Y(N560) );
  AOI21X1TF U544 ( .A0(N119), .A1(N651), .B0(N976), .Y(N562) );
  INVX2TF U545 ( .A(SUM_AB[0]), .Y(N976) );
  AOI32X1TF U546 ( .A0(N461), .A1(N460), .A2(N459), .B0(N475), .B1(N154), .Y(
        N712) );
  OAI211X1TF U547 ( .A0(N507), .A1(N997), .B0(N456), .C0(N455), .Y(N457) );
  AOI22X1TF U548 ( .A0(DIVISION_HEAD[12]), .A1(N95), .B0(X_IN[12]), .B1(N102), 
        .Y(N455) );
  AOI22X1TF U549 ( .A0(DIVISION_HEAD[11]), .A1(N806), .B0(DIVISION_HEAD[10]), 
        .B1(N131), .Y(N456) );
  OAI22X1TF U550 ( .A0(N463), .A1(N609), .B0(N559), .B1(N498), .Y(N458) );
  OAI22X1TF U551 ( .A0(N196), .A1(N753), .B0(N761), .B1(N177), .Y(N688) );
  AOI211X1TF U552 ( .A0(N992), .A1(N797), .B0(N752), .C0(N751), .Y(N753) );
  OAI211X1TF U553 ( .A0(N750), .A1(N749), .B0(N757), .C0(N748), .Y(N751) );
  AOI22X1TF U554 ( .A0(DIVISION_REMA[7]), .A1(N120), .B0(SUM_AB[6]), .B1(N145), 
        .Y(N748) );
  OAI21X1TF U555 ( .A0(N206), .A1(N100), .B0(N746), .Y(N752) );
  AOI22X1TF U556 ( .A0(Y_IN[6]), .A1(N791), .B0(DIVISION_REMA[5]), .B1(N736), 
        .Y(N746) );
  AOI21X1TF U557 ( .A0(SUM_AB[6]), .A1(N443), .B0(N453), .Y(N992) );
  OAI22X1TF U558 ( .A0(N513), .A1(N362), .B0(N361), .B1(N179), .Y(N723) );
  AOI211X1TF U559 ( .A0(N493), .A1(N1013), .B0(N359), .C0(N358), .Y(N362) );
  OAI31X1TF U560 ( .A0(XTEMP[12]), .A1(N360), .A2(N509), .B0(N357), .Y(N358)
         );
  AOI22X1TF U561 ( .A0(XTEMP[11]), .A1(N131), .B0(N139), .B1(N444), .Y(N357)
         );
  INVX2TF U562 ( .A(INTADD_0_N1), .Y(N464) );
  OAI22X1TF U563 ( .A0(N119), .A1(N1018), .B0(N502), .B1(N100), .Y(N359) );
  OAI21X1TF U564 ( .A0(N814), .A1(N556), .B0(N555), .Y(N706) );
  OAI21X1TF U565 ( .A0(N814), .A1(N806), .B0(DIVISION_HEAD[3]), .Y(N555) );
  AOI211X1TF U566 ( .A0(DIVISION_HEAD[2]), .A1(N131), .B0(N554), .C0(N553), 
        .Y(N556) );
  AOI22X1TF U567 ( .A0(N800), .A1(SUM_AB[3]), .B0(N1013), .B1(N797), .Y(N550)
         );
  NOR2X1TF U568 ( .A(N1018), .B(N1014), .Y(N1013) );
  AOI22X1TF U569 ( .A0(N941), .A1(SUM_AB[12]), .B0(N106), .B1(N137), .Y(N551)
         );
  OAI22X1TF U570 ( .A0(N549), .A1(N804), .B0(N548), .B1(N100), .Y(N554) );
  OAI22X1TF U571 ( .A0(N196), .A1(N655), .B0(N761), .B1(N184), .Y(N693) );
  AOI21X1TF U572 ( .A0(SUM_AB[1]), .A1(N146), .B0(N654), .Y(N655) );
  AOI22X1TF U573 ( .A0(DIVISION_REMA[0]), .A1(N736), .B0(N797), .B1(N977), .Y(
        N652) );
  AOI21X1TF U574 ( .A0(SUM_AB[1]), .A1(SUM_AB[0]), .B0(N403), .Y(N977) );
  AOI22X1TF U575 ( .A0(Y_IN[1]), .A1(N791), .B0(DIVISION_REMA[2]), .B1(N125), 
        .Y(N653) );
  AOI22X1TF U576 ( .A0(N196), .A1(N149), .B0(N781), .B1(N780), .Y(N686) );
  AOI211X1TF U577 ( .A0(DIVISION_REMA[7]), .A1(N736), .B0(N779), .C0(N778), 
        .Y(N781) );
  OAI211X1TF U578 ( .A0(N174), .A1(N777), .B0(N776), .C0(N775), .Y(N778) );
  AOI22X1TF U579 ( .A0(N774), .A1(N773), .B0(N998), .B1(N797), .Y(N775) );
  AOI21X1TF U580 ( .A0(SUM_AB[8]), .A1(N462), .B0(N477), .Y(N998) );
  AOI32X1TF U581 ( .A0(N772), .A1(N771), .A2(N770), .B0(N769), .B1(N771), .Y(
        N773) );
  AOI22X1TF U582 ( .A0(DIVISION_REMA[8]), .A1(N763), .B0(SUM_AB[8]), .B1(N145), 
        .Y(N776) );
  AOI22X1TF U583 ( .A0(N475), .A1(N156), .B0(N441), .B1(N460), .Y(N714) );
  AOI21X1TF U584 ( .A0(DIVISION_HEAD[8]), .A1(N131), .B0(N434), .Y(N435) );
  OAI22X1TF U585 ( .A0(N156), .A1(N454), .B0(N507), .B1(N991), .Y(N434) );
  AOI22X1TF U586 ( .A0(DIVISION_HEAD[10]), .A1(N95), .B0(X_IN[10]), .B1(N101), 
        .Y(N437) );
  OAI22X1TF U587 ( .A0(N442), .A1(N609), .B0(N559), .B1(N476), .Y(N440) );
  OAI22X1TF U588 ( .A0(N196), .A1(N741), .B0(N761), .B1(N176), .Y(N690) );
  AOI211X1TF U589 ( .A0(SUM_AB[4]), .A1(N146), .B0(N740), .C0(N739), .Y(N741)
         );
  OAI211X1TF U590 ( .A0(N738), .A1(N100), .B0(N757), .C0(N737), .Y(N739) );
  AOI22X1TF U591 ( .A0(DIVISION_REMA[5]), .A1(N125), .B0(N797), .B1(N986), .Y(
        N737) );
  AOI21X1TF U592 ( .A0(SUM_AB[4]), .A1(N422), .B0(N433), .Y(N986) );
  OAI22X1TF U593 ( .A0(N206), .A1(N804), .B0(N171), .B1(N98), .Y(N740) );
  OAI22X1TF U594 ( .A0(N196), .A1(N730), .B0(N761), .B1(N150), .Y(N692) );
  AOI211X1TF U595 ( .A0(SUM_AB[2]), .A1(N146), .B0(N729), .C0(N728), .Y(N730)
         );
  OAI211X1TF U596 ( .A0(N727), .A1(N100), .B0(N757), .C0(N656), .Y(N728) );
  AOI22X1TF U597 ( .A0(DIVISION_REMA[3]), .A1(N125), .B0(N797), .B1(N980), .Y(
        N656) );
  AOI21X1TF U598 ( .A0(SUM_AB[2]), .A1(N404), .B0(N414), .Y(N980) );
  NOR2X1TF U599 ( .A(SUM_AB[0]), .B(SUM_AB[1]), .Y(N403) );
  OAI22X1TF U600 ( .A0(N738), .A1(N804), .B0(N184), .B1(N98), .Y(N729) );
  AOI32X1TF U601 ( .A0(N421), .A1(N460), .A2(N420), .B0(N475), .B1(N423), .Y(
        N716) );
  AOI211X1TF U602 ( .A0(DIVISION_HEAD[8]), .A1(N96), .B0(N419), .C0(N418), .Y(
        N420) );
  OAI211X1TF U603 ( .A0(N559), .A1(N452), .B0(N417), .C0(N416), .Y(N418) );
  AOI21X1TF U604 ( .A0(DIVISION_HEAD[6]), .A1(N736), .B0(N415), .Y(N416) );
  OAI22X1TF U605 ( .A0(N423), .A1(N454), .B0(N507), .B1(N985), .Y(N415) );
  INVX2TF U606 ( .A(N493), .Y(N507) );
  NOR2X2TF U607 ( .A(N393), .B(N1018), .Y(N493) );
  INVX2TF U608 ( .A(N609), .Y(N444) );
  NAND2X2TF U609 ( .A(MODE_TYPE[1]), .B(N356), .Y(N609) );
  OAI21X1TF U610 ( .A0(N502), .A1(N749), .B0(N412), .Y(N419) );
  AOI22X1TF U611 ( .A0(X_IN[8]), .A1(N102), .B0(N82), .B1(N137), .Y(N412) );
  INVX2TF U612 ( .A(N807), .Y(N749) );
  AOI31X1TF U613 ( .A0(N941), .A1(N73), .A2(N564), .B0(N353), .Y(N384) );
  OAI211X1TF U614 ( .A0(N73), .A1(N378), .B0(N363), .C0(N352), .Y(N353) );
  OAI211X1TF U615 ( .A0(N960), .A1(N351), .B0(N567), .C0(N601), .Y(N352) );
  NOR2X1TF U616 ( .A(N375), .B(N944), .Y(N363) );
  INVX2TF U617 ( .A(N393), .Y(N375) );
  INVX2TF U618 ( .A(N618), .Y(N378) );
  NOR2X1TF U619 ( .A(N158), .B(N750), .Y(INTADD_0_CI) );
  INVX2TF U620 ( .A(X_IN[0]), .Y(N750) );
  NOR2X1TF U621 ( .A(PRE_WORK), .B(N368), .Y(N603) );
  INVX2TF U622 ( .A(N600), .Y(N567) );
  OAI211X1TF U623 ( .A0(N862), .A1(N861), .B0(N860), .C0(N859), .Y(N678) );
  AOI32X1TF U624 ( .A0(N937), .A1(OPER_B[4]), .A2(N858), .B0(N890), .B1(
        OPER_B[4]), .Y(N859) );
  AOI211X1TF U625 ( .A0(N864), .A1(OPER_B[5]), .B0(N857), .C0(N856), .Y(N860)
         );
  OAI31X1TF U626 ( .A0(N934), .A1(OPER_A[4]), .A2(N855), .B0(N210), .Y(N856)
         );
  AOI21X1TF U627 ( .A0(N113), .A1(C152_DATA4_4), .B0(N211), .Y(N210) );
  NOR3X1TF U628 ( .A(OPER_B[4]), .B(N858), .C(N116), .Y(N857) );
  AOI21X1TF U629 ( .A0(N931), .A1(N855), .B0(N854), .Y(N861) );
  OAI211X1TF U630 ( .A0(N830), .A1(N832), .B0(N829), .C0(N212), .Y(N681) );
  AOI211X1TF U631 ( .A0(N114), .A1(C152_DATA4_1), .B0(N826), .C0(N891), .Y(
        N212) );
  OAI31X1TF U632 ( .A0(OPER_B[1]), .A1(N116), .A2(N189), .B0(N825), .Y(N826)
         );
  AOI211X1TF U633 ( .A0(N864), .A1(OPER_B[2]), .B0(N828), .C0(N827), .Y(N829)
         );
  NOR3X1TF U634 ( .A(N831), .B(OPER_A[1]), .C(N934), .Y(N827) );
  OAI32X1TF U635 ( .A0(N187), .A1(OPER_B[0]), .A2(N116), .B0(N935), .B1(N187), 
        .Y(N828) );
  AOI21X1TF U636 ( .A0(N931), .A1(N831), .B0(N854), .Y(N830) );
  INVX2TF U637 ( .A(N932), .Y(N854) );
  NOR2X1TF U638 ( .A(N104), .B(N159), .Y(FOUT[11]) );
  AOI211X1TF U639 ( .A0(N114), .A1(C152_DATA4_5), .B0(N866), .C0(N215), .Y(
        N216) );
  OAI31X1TF U640 ( .A0(OPER_B[5]), .A1(N865), .A2(N116), .B0(N905), .Y(N866)
         );
  OAI211X1TF U641 ( .A0(SIGN_Y), .A1(N965), .B0(N225), .C0(N972), .Y(N905) );
  AOI22X1TF U642 ( .A0(N864), .A1(OPER_B[6]), .B0(N863), .B1(N868), .Y(N873)
         );
  NOR2X1TF U643 ( .A(N934), .B(OPER_A[5]), .Y(N863) );
  INVX2TF U644 ( .A(N894), .Y(N864) );
  AOI22X1TF U645 ( .A0(OPER_B[5]), .A1(N870), .B0(OPER_A[5]), .B1(N869), .Y(
        N872) );
  OAI21X1TF U646 ( .A0(N934), .A1(N868), .B0(N932), .Y(N869) );
  OAI21X1TF U647 ( .A0(N116), .A1(N867), .B0(N935), .Y(N870) );
  OR2X2TF U648 ( .A(N930), .B(N891), .Y(N211) );
  NOR2X1TF U649 ( .A(N967), .B(N836), .Y(N876) );
  INVX2TF U650 ( .A(N935), .Y(N890) );
  NOR3X1TF U651 ( .A(N73), .B(N182), .C(N965), .Y(N964) );
  OAI22X1TF U652 ( .A0(N133), .A1(N206), .B0(OFFSET[2]), .B1(N207), .Y(C2_Z_4)
         );
  INVX2TF U653 ( .A(Y_IN[4]), .Y(N206) );
  OAI22X1TF U654 ( .A0(N133), .A1(N205), .B0(OFFSET[3]), .B1(N207), .Y(C2_Z_5)
         );
  OAI22X1TF U655 ( .A0(N132), .A1(N204), .B0(OFFSET[4]), .B1(N207), .Y(C2_Z_6)
         );
  OAI22X1TF U656 ( .A0(N132), .A1(N198), .B0(OFFSET[5]), .B1(N207), .Y(C2_Z_7)
         );
  NOR2X1TF U657 ( .A(OPER_B[9]), .B(N908), .Y(N923) );
  NOR2X1TF U658 ( .A(N875), .B(OPER_B[6]), .Y(N892) );
  INVX2TF U659 ( .A(N879), .Y(N875) );
  NOR2X1TF U660 ( .A(OPER_B[5]), .B(N867), .Y(N879) );
  NOR2X1TF U661 ( .A(OPER_B[3]), .B(N847), .Y(N858) );
  AOI211X1TF U662 ( .A0(N61), .A1(N965), .B0(SIGN_Y), .C0(N910), .Y(N930) );
  NOR2X1TF U663 ( .A(OPER_A[9]), .B(N909), .Y(N917) );
  NOR2X1TF U664 ( .A(OPER_A[7]), .B(N893), .Y(N898) );
  NOR2X1TF U665 ( .A(OPER_A[5]), .B(N868), .Y(N882) );
  NOR2X1TF U666 ( .A(OPER_A[3]), .B(N846), .Y(N855) );
  OAI211X1TF U667 ( .A0(N181), .A1(N938), .B0(N853), .C0(N852), .Y(N679) );
  AOI211X1TF U668 ( .A0(OPER_A[3]), .A1(N851), .B0(N850), .C0(N849), .Y(N852)
         );
  OAI31X1TF U669 ( .A0(N934), .A1(OPER_A[3]), .A2(N848), .B0(N209), .Y(N849)
         );
  AOI21X1TF U670 ( .A0(C152_DATA4_3), .A1(N113), .B0(N906), .Y(N209) );
  NOR2X1TF U671 ( .A(N61), .B(N910), .Y(N906) );
  OAI21X1TF U672 ( .A0(N133), .A1(N317), .B0(N207), .Y(C2_Z_1) );
  OAI22X1TF U673 ( .A0(N133), .A1(N731), .B0(OFFSET[1]), .B1(N207), .Y(C2_Z_3)
         );
  OAI32X1TF U674 ( .A0(N188), .A1(N115), .A2(N847), .B0(N935), .B1(N188), .Y(
        N850) );
  INVX2TF U675 ( .A(N874), .Y(N921) );
  AOI32X1TF U676 ( .A0(N606), .A1(N350), .A2(N824), .B0(N946), .B1(N349), .Y(
        N874) );
  INVX2TF U677 ( .A(N940), .Y(N946) );
  OAI21X1TF U678 ( .A0(N934), .A1(N846), .B0(N932), .Y(N851) );
  INVX2TF U679 ( .A(N837), .Y(N912) );
  AOI21X1TF U680 ( .A0(N565), .A1(N349), .B0(N564), .Y(N837) );
  INVX2TF U681 ( .A(N848), .Y(N846) );
  NOR3X1TF U682 ( .A(OPER_A[2]), .B(OPER_A[1]), .C(OPER_A[0]), .Y(N848) );
  INVX2TF U683 ( .A(N931), .Y(N934) );
  NOR2X2TF U684 ( .A(N924), .B(N916), .Y(N931) );
  INVX2TF U685 ( .A(N904), .Y(N924) );
  AOI31X1TF U686 ( .A0(N937), .A1(N188), .A2(N847), .B0(N888), .Y(N853) );
  OAI21X1TF U687 ( .A0(N975), .A1(N910), .B0(N843), .Y(N888) );
  INVX2TF U688 ( .A(N910), .Y(N225) );
  INVX2TF U689 ( .A(N348), .Y(N959) );
  INVX2TF U690 ( .A(N566), .Y(N949) );
  NOR2X1TF U691 ( .A(OPER_B[1]), .B(OPER_B[0]), .Y(N839) );
  INVX2TF U692 ( .A(N349), .Y(N350) );
  INVX2TF U693 ( .A(N606), .Y(N823) );
  NOR2X2TF U694 ( .A(N604), .B(N632), .Y(N824) );
  AOI221X1TF U695 ( .A0(N128), .A1(N164), .B0(N186), .B1(N91), .C0(N819), .Y(
        N820) );
  AOI22X1TF U696 ( .A0(\INDEX[2] ), .A1(N90), .B0(N124), .B1(\RSHT_BITS[3] ), 
        .Y(N818) );
  AOI32X1TF U697 ( .A0(N940), .A1(N953), .A2(N372), .B0(N955), .B1(N953), .Y(
        N346) );
  OR2X2TF U698 ( .A(N632), .B(N152), .Y(N372) );
  INVX2TF U699 ( .A(N604), .Y(N643) );
  OAI21X1TF U700 ( .A0(N348), .A1(N939), .B0(N344), .Y(N608) );
  OAI21X1TF U701 ( .A0(N571), .A1(N565), .B0(N345), .Y(N344) );
  NOR2X2TF U702 ( .A(\RSHT_BITS[3] ), .B(N592), .Y(N606) );
  NOR3X1TF U703 ( .A(N121), .B(N122), .C(N954), .Y(N822) );
  INVX2TF U704 ( .A(N960), .Y(N967) );
  NOR2X1TF U705 ( .A(SIGN_Y), .B(N117), .Y(N907) );
  OAI22X1TF U706 ( .A0(Y_IN[12]), .A1(N178), .B0(N340), .B1(N339), .Y(N341) );
  OAI31X1TF U707 ( .A0(N338), .A1(DIVISION_HEAD[10]), .A2(N548), .B0(N337), 
        .Y(N339) );
  AOI22X1TF U708 ( .A0(Y_IN[11]), .A1(N154), .B0(N336), .B1(N335), .Y(N337) );
  OAI22X1TF U709 ( .A0(DIVISION_HEAD[8]), .A1(N762), .B0(DIVISION_HEAD[9]), 
        .B1(N784), .Y(N335) );
  INVX2TF U710 ( .A(N334), .Y(N336) );
  NOR2X1TF U711 ( .A(Y_IN[11]), .B(N154), .Y(N338) );
  AOI211X1TF U712 ( .A0(DIVISION_HEAD[8]), .A1(N762), .B0(N333), .C0(N334), 
        .Y(N340) );
  OAI21X1TF U713 ( .A0(Y_IN[11]), .A1(N154), .B0(N332), .Y(N334) );
  AOI22X1TF U714 ( .A0(DIVISION_HEAD[10]), .A1(N548), .B0(DIVISION_HEAD[9]), 
        .B1(N784), .Y(N332) );
  AOI21X1TF U715 ( .A0(N89), .A1(N423), .B0(N331), .Y(N333) );
  AOI211X1TF U716 ( .A0(N330), .A1(DIVISION_HEAD[6]), .B0(N329), .C0(N328), 
        .Y(N331) );
  NOR2X1TF U717 ( .A(N89), .B(N423), .Y(N329) );
  AOI211X1TF U718 ( .A0(N326), .A1(DIVISION_HEAD[4]), .B0(N325), .C0(N324), 
        .Y(N327) );
  NOR2X1TF U719 ( .A(Y_IN[5]), .B(N514), .Y(N325) );
  AOI21X1TF U720 ( .A0(Y_IN[3]), .A1(N649), .B0(N323), .Y(N326) );
  OAI32X1TF U721 ( .A0(N322), .A1(DIVISION_HEAD[2]), .A2(N738), .B0(N321), 
        .B1(N322), .Y(N323) );
  OAI211X1TF U722 ( .A0(Y_IN[2]), .A1(N168), .B0(N320), .C0(N319), .Y(N321) );
  NOR2X1TF U723 ( .A(Y_IN[3]), .B(N649), .Y(N322) );
  INVX2TF U724 ( .A(Y_IN[12]), .Y(N549) );
  OAI21X1TF U725 ( .A0(N154), .A1(N104), .B0(N241), .Y(FOUT[7]) );
  AOI21X1TF U726 ( .A0(N224), .A1(DIVISION_REMA[7]), .B0(N240), .Y(N241) );
  OAI22X1TF U727 ( .A0(N174), .A1(N86), .B0(N529), .B1(N83), .Y(N240) );
  OAI21X1TF U728 ( .A0(N160), .A1(N104), .B0(N239), .Y(FOUT[6]) );
  AOI21X1TF U729 ( .A0(N224), .A1(DIVISION_REMA[6]), .B0(N238), .Y(N239) );
  OAI22X1TF U730 ( .A0(N178), .A1(N84), .B0(N149), .B1(N86), .Y(N238) );
  OAI21X1TF U731 ( .A0(N761), .A1(N173), .B0(N760), .Y(N687) );
  OAI21X1TF U732 ( .A0(N759), .A1(N758), .B0(N780), .Y(N760) );
  INVX2TF U733 ( .A(N196), .Y(N780) );
  OAI211X1TF U734 ( .A0(N149), .A1(N777), .B0(N757), .C0(N756), .Y(N758) );
  AOI22X1TF U735 ( .A0(DIVISION_REMA[6]), .A1(N736), .B0(SUM_AB[7]), .B1(N145), 
        .Y(N756) );
  OAI211X1TF U736 ( .A0(N810), .A1(N997), .B0(N755), .C0(N754), .Y(N759) );
  OAI21X1TF U737 ( .A0(N453), .A1(N452), .B0(N462), .Y(N997) );
  NOR2X1TF U738 ( .A(N104), .B(N179), .Y(FOUT[12]) );
  OAI22X1TF U739 ( .A0(N196), .A1(N745), .B0(N761), .B1(N172), .Y(N689) );
  AOI211X1TF U740 ( .A0(SUM_AB[5]), .A1(N146), .B0(N744), .C0(N743), .Y(N745)
         );
  OAI211X1TF U741 ( .A0(N810), .A1(N991), .B0(N757), .C0(N742), .Y(N743) );
  OAI21X1TF U742 ( .A0(N433), .A1(N432), .B0(N443), .Y(N991) );
  INVX2TF U743 ( .A(N804), .Y(N791) );
  OAI22X1TF U744 ( .A0(N196), .A1(N735), .B0(N761), .B1(N171), .Y(N691) );
  AOI211X1TF U745 ( .A0(SUM_AB[3]), .A1(N146), .B0(N734), .C0(N733), .Y(N735)
         );
  OAI211X1TF U746 ( .A0(N810), .A1(N985), .B0(N757), .C0(N732), .Y(N733) );
  AOI222X4TF U747 ( .A0(N767), .A1(N101), .B0(N765), .B1(N136), .C0(N558), 
        .C1(N807), .Y(N757) );
  OAI21X1TF U748 ( .A0(N414), .A1(N413), .B0(N422), .Y(N985) );
  OAI22X1TF U749 ( .A0(N731), .A1(N804), .B0(N150), .B1(N98), .Y(N734) );
  NOR3X1TF U750 ( .A(N774), .B(N131), .C(N557), .Y(N782) );
  AOI32X1TF U751 ( .A0(N790), .A1(N816), .A2(N789), .B0(N814), .B1(N174), .Y(
        N685) );
  OAI211X1TF U752 ( .A0(N810), .A1(N1003), .B0(N786), .C0(N785), .Y(N787) );
  AOI22X1TF U753 ( .A0(DIVISION_HEAD[1]), .A1(N125), .B0(X_IN[1]), .B1(N101), 
        .Y(N785) );
  OAI21X1TF U754 ( .A0(N477), .A1(N476), .B0(N486), .Y(N1003) );
  OAI21X1TF U755 ( .A0(N784), .A1(N804), .B0(N783), .Y(N788) );
  AOI22X1TF U756 ( .A0(DIVISION_REMA[8]), .A1(N131), .B0(N800), .B1(SUM_AB[0]), 
        .Y(N783) );
  AOI22X1TF U757 ( .A0(DIVISION_HEAD[0]), .A1(N806), .B0(SUM_AB[9]), .B1(N146), 
        .Y(N790) );
  OAI21X1TF U758 ( .A0(N156), .A1(N103), .B0(N237), .Y(FOUT[5]) );
  AOI21X1TF U759 ( .A0(N224), .A1(DIVISION_REMA[5]), .B0(N236), .Y(N237) );
  OAI22X1TF U760 ( .A0(N154), .A1(N83), .B0(N173), .B1(N85), .Y(N236) );
  AOI32X1TF U761 ( .A0(N817), .A1(N816), .A2(N815), .B0(N814), .B1(N168), .Y(
        N683) );
  AOI211X1TF U762 ( .A0(DIVISION_HEAD[3]), .A1(N125), .B0(N812), .C0(N811), 
        .Y(N815) );
  OAI211X1TF U763 ( .A0(N810), .A1(N1009), .B0(N809), .C0(N808), .Y(N811) );
  AND2X2TF U764 ( .A(N764), .B(N769), .Y(N766) );
  INVX2TF U765 ( .A(N385), .Y(N774) );
  AOI22X1TF U766 ( .A0(DIVISION_HEAD[1]), .A1(N131), .B0(DIVISION_HEAD[2]), 
        .B1(N806), .Y(N809) );
  INVX2TF U767 ( .A(N454), .Y(N806) );
  OAI21X1TF U768 ( .A0(N499), .A1(N498), .B0(N1014), .Y(N1009) );
  INVX2TF U769 ( .A(SUM_AB[11]), .Y(N498) );
  INVX2TF U770 ( .A(SUM_AB[9]), .Y(N476) );
  INVX2TF U771 ( .A(SUM_AB[7]), .Y(N452) );
  NOR2X1TF U772 ( .A(SUM_AB[6]), .B(N443), .Y(N453) );
  INVX2TF U773 ( .A(SUM_AB[5]), .Y(N432) );
  NOR2X1TF U774 ( .A(SUM_AB[4]), .B(N422), .Y(N433) );
  INVX2TF U775 ( .A(SUM_AB[3]), .Y(N413) );
  NOR3X1TF U776 ( .A(SUM_AB[0]), .B(SUM_AB[2]), .C(SUM_AB[1]), .Y(N414) );
  INVX2TF U777 ( .A(N797), .Y(N810) );
  NOR2X2TF U778 ( .A(N1018), .B(N651), .Y(N797) );
  INVX2TF U779 ( .A(SUM_AB[12]), .Y(N1018) );
  OAI21X1TF U780 ( .A0(N805), .A1(N804), .B0(N803), .Y(N812) );
  INVX2TF U781 ( .A(N99), .Y(N802) );
  NAND2X2TF U782 ( .A(N356), .B(N315), .Y(N804) );
  INVX2TF U783 ( .A(N814), .Y(N816) );
  INVX2TF U784 ( .A(N356), .Y(N640) );
  AOI31X1TF U785 ( .A0(N122), .A1(N383), .A2(N382), .B0(N381), .Y(N547) );
  INVX2TF U786 ( .A(N308), .Y(N765) );
  OAI211X1TF U787 ( .A0(X_IN[12]), .A1(N548), .B0(N307), .C0(N306), .Y(N308)
         );
  OAI22X1TF U788 ( .A0(Y_IN[10]), .A1(N305), .B0(N304), .B1(N303), .Y(N306) );
  OAI22X1TF U789 ( .A0(X_IN[10]), .A1(N302), .B0(N138), .B1(N784), .Y(N303) );
  OAI21X1TF U790 ( .A0(Y_IN[9]), .A1(N201), .B0(Y_IN[8]), .Y(N302) );
  AOI211X1TF U791 ( .A0(X_IN[10]), .A1(N762), .B0(N301), .C0(N300), .Y(N304)
         );
  AOI21X1TF U792 ( .A0(N89), .A1(N500), .B0(N299), .Y(N300) );
  AOI211X1TF U793 ( .A0(X_IN[8]), .A1(N298), .B0(N297), .C0(N296), .Y(N299) );
  NOR2X1TF U794 ( .A(N89), .B(N500), .Y(N297) );
  AOI21X1TF U795 ( .A0(N197), .A1(N468), .B0(N295), .Y(N298) );
  AOI211X1TF U796 ( .A0(X_IN[6]), .A1(N294), .B0(N293), .C0(N292), .Y(N295) );
  NOR2X1TF U797 ( .A(N197), .B(N468), .Y(N293) );
  AOI32X1TF U798 ( .A0(N291), .A1(N290), .A2(N319), .B0(N289), .B1(N290), .Y(
        N294) );
  OAI22X1TF U799 ( .A0(X_IN[4]), .A1(N738), .B0(N106), .B1(N731), .Y(N289) );
  OAI32X1TF U800 ( .A0(N288), .A1(N93), .A2(N317), .B0(X_IN[2]), .B1(N288), 
        .Y(N291) );
  INVX2TF U801 ( .A(X_IN[7]), .Y(N468) );
  INVX2TF U802 ( .A(X_IN[9]), .Y(N500) );
  NOR2X1TF U803 ( .A(Y_IN[9]), .B(N201), .Y(N301) );
  NOR2X1TF U804 ( .A(Y_IN[12]), .B(Y_IN[11]), .Y(N307) );
  INVX2TF U805 ( .A(N770), .Y(N558) );
  OR2X2TF U806 ( .A(MODE_TYPE[0]), .B(N315), .Y(N769) );
  INVX2TF U807 ( .A(MODE_TYPE[1]), .Y(N315) );
  OAI31X1TF U808 ( .A0(N286), .A1(N139), .A2(N548), .B0(N285), .Y(N287) );
  OAI31X1TF U809 ( .A0(N284), .A1(N283), .A2(N282), .B0(N281), .Y(N285) );
  AOI22X1TF U810 ( .A0(N138), .A1(N548), .B0(X_IN[12]), .B1(N805), .Y(N281) );
  INVX2TF U811 ( .A(Y_IN[11]), .Y(N805) );
  NOR2X1TF U812 ( .A(X_IN[10]), .B(N784), .Y(N282) );
  AOI211X1TF U813 ( .A0(X_IN[10]), .A1(N784), .B0(X_IN[9]), .C0(N762), .Y(N283) );
  INVX2TF U814 ( .A(Y_IN[9]), .Y(N784) );
  AOI211X1TF U815 ( .A0(X_IN[9]), .A1(N762), .B0(N280), .C0(N279), .Y(N284) );
  AOI21X1TF U816 ( .A0(N89), .A1(N488), .B0(N278), .Y(N279) );
  AOI211X1TF U817 ( .A0(N277), .A1(X_IN[7]), .B0(N276), .C0(N275), .Y(N278) );
  NOR2X1TF U818 ( .A(N89), .B(N488), .Y(N276) );
  AOI21X1TF U819 ( .A0(N197), .A1(N463), .B0(N274), .Y(N277) );
  AOI211X1TF U820 ( .A0(N273), .A1(N106), .B0(N272), .C0(N271), .Y(N274) );
  NOR2X1TF U821 ( .A(N197), .B(N463), .Y(N272) );
  AOI211X1TF U822 ( .A0(Y_IN[3]), .A1(N442), .B0(N270), .C0(N269), .Y(N273) );
  AOI211X1TF U823 ( .A0(X_IN[4]), .A1(N731), .B0(N94), .C0(N738), .Y(N269) );
  INVX2TF U824 ( .A(Y_IN[3]), .Y(N731) );
  OAI32X1TF U825 ( .A0(N268), .A1(X_IN[2]), .A2(N317), .B0(X_IN[1]), .B1(N268), 
        .Y(N270) );
  OAI211X1TF U826 ( .A0(Y_IN[3]), .A1(N442), .B0(N267), .C0(N319), .Y(N268) );
  INVX2TF U827 ( .A(Y_IN[0]), .Y(N727) );
  INVX2TF U828 ( .A(Y_IN[1]), .Y(N317) );
  AOI22X1TF U829 ( .A0(N93), .A1(N738), .B0(X_IN[2]), .B1(N318), .Y(N267) );
  INVX2TF U830 ( .A(Y_IN[2]), .Y(N738) );
  INVX2TF U831 ( .A(X_IN[4]), .Y(N442) );
  INVX2TF U832 ( .A(X_IN[6]), .Y(N463) );
  INVX2TF U833 ( .A(X_IN[8]), .Y(N488) );
  NOR2X1TF U834 ( .A(Y_IN[9]), .B(N502), .Y(N280) );
  INVX2TF U835 ( .A(X_IN[10]), .Y(N502) );
  INVX2TF U836 ( .A(Y_IN[8]), .Y(N762) );
  INVX2TF U837 ( .A(Y_IN[10]), .Y(N548) );
  NOR2X1TF U838 ( .A(Y_IN[11]), .B(N305), .Y(N286) );
  INVX2TF U839 ( .A(X_IN[12]), .Y(N305) );
  INVX2TF U840 ( .A(N342), .Y(N383) );
  AOI22X1TF U841 ( .A0(N800), .A1(SUM_AB[2]), .B0(SUM_AB[11]), .B1(N146), .Y(
        N817) );
  INVX2TF U842 ( .A(N312), .Y(N628) );
  OAI21X1TF U843 ( .A0(N179), .A1(N112), .B0(N260), .Y(OPER_A[12]) );
  OAI21X1TF U844 ( .A0(N423), .A1(N111), .B0(N250), .Y(OPER_A[3]) );
  OAI21X1TF U845 ( .A0(N155), .A1(N112), .B0(N251), .Y(OPER_A[4]) );
  OAI21X1TF U846 ( .A0(N156), .A1(N112), .B0(N252), .Y(OPER_A[5]) );
  OAI21X1TF U847 ( .A0(N160), .A1(N112), .B0(N253), .Y(OPER_A[6]) );
  OAI21X1TF U848 ( .A0(N154), .A1(N112), .B0(N254), .Y(OPER_A[7]) );
  OAI21X1TF U849 ( .A0(N178), .A1(N112), .B0(N255), .Y(OPER_A[8]) );
  OAI21X1TF U850 ( .A0(N112), .A1(N529), .B0(N256), .Y(OPER_A[9]) );
  OAI21X1TF U851 ( .A0(N112), .A1(N161), .B0(N257), .Y(OPER_A[10]) );
  OAI21X1TF U852 ( .A0(N112), .A1(N159), .B0(N258), .Y(OPER_A[11]) );
  OAI21X1TF U853 ( .A0(N157), .A1(N111), .B0(N249), .Y(OPER_A[2]) );
  INVX2TF U854 ( .A(N559), .Y(N800) );
  OAI21X1TF U855 ( .A0(N514), .A1(N103), .B0(N229), .Y(FOUT[1]) );
  AOI21X1TF U856 ( .A0(N224), .A1(DIVISION_REMA[1]), .B0(N228), .Y(N229) );
  OAI22X1TF U857 ( .A0(N423), .A1(N83), .B0(N171), .B1(N85), .Y(N228) );
  NOR2X1TF U858 ( .A(N342), .B(N373), .Y(ALU_IS_DONE) );
  OAI211X1TF U859 ( .A0(N157), .A1(N84), .B0(N227), .C0(N226), .Y(FOUT[0]) );
  OAI21X1TF U860 ( .A0(N178), .A1(N104), .B0(N243), .Y(FOUT[8]) );
  AOI21X1TF U861 ( .A0(N224), .A1(DIVISION_REMA[8]), .B0(N242), .Y(N243) );
  OAI22X1TF U862 ( .A0(N175), .A1(N86), .B0(N161), .B1(N84), .Y(N242) );
  OAI21X1TF U863 ( .A0(N155), .A1(N103), .B0(N235), .Y(FOUT[4]) );
  AOI21X1TF U864 ( .A0(N224), .A1(DIVISION_REMA[4]), .B0(N234), .Y(N235) );
  OAI22X1TF U865 ( .A0(N160), .A1(N84), .B0(N177), .B1(N86), .Y(N234) );
  OAI21X1TF U866 ( .A0(N423), .A1(N103), .B0(N233), .Y(FOUT[3]) );
  AOI21X1TF U867 ( .A0(N224), .A1(DIVISION_REMA[3]), .B0(N232), .Y(N233) );
  OAI22X1TF U868 ( .A0(N156), .A1(N84), .B0(N172), .B1(N85), .Y(N232) );
  OAI21X1TF U869 ( .A0(N157), .A1(N103), .B0(N231), .Y(FOUT[2]) );
  AOI21X1TF U870 ( .A0(N224), .A1(DIVISION_REMA[2]), .B0(N230), .Y(N231) );
  OAI22X1TF U871 ( .A0(N155), .A1(N83), .B0(N176), .B1(N85), .Y(N230) );
  AOI21X1TF U872 ( .A0(N127), .A1(N472), .B0(N471), .Y(N473) );
  AOI22X1TF U873 ( .A0(N126), .A1(N465), .B0(SUM_AB[8]), .B1(N134), .Y(N467)
         );
  AOI22X1TF U874 ( .A0(N127), .A1(\INTADD_0_SUM[5] ), .B0(N800), .B1(
        SUM_AB[10]), .Y(N448) );
  AOI22X1TF U875 ( .A0(N127), .A1(\INTADD_0_SUM[3] ), .B0(SUM_AB[4]), .B1(N135), .Y(N431) );
  AOI31X1TF U876 ( .A0(X_IN[0]), .A1(N127), .A2(N158), .B0(N389), .Y(N390) );
  AOI22X1TF U877 ( .A0(N127), .A1(\INTADD_0_SUM[0] ), .B0(SUM_AB[1]), .B1(N135), .Y(N401) );
  AOI31X1TF U878 ( .A0(N126), .A1(N161), .A2(N494), .B0(N489), .Y(N490) );
  AOI22X1TF U879 ( .A0(N127), .A1(\INTADD_0_SUM[1] ), .B0(SUM_AB[2]), .B1(N135), .Y(N411) );
  AOI31X1TF U880 ( .A0(N127), .A1(N159), .A2(N510), .B0(N508), .Y(N512) );
  AOI22X1TF U881 ( .A0(N127), .A1(\INTADD_0_SUM[6] ), .B0(SUM_AB[7]), .B1(N135), .Y(N461) );
  AOI21X1TF U882 ( .A0(N127), .A1(N360), .B0(N513), .Y(N361) );
  AOI22X1TF U883 ( .A0(N126), .A1(\INTADD_0_SUM[4] ), .B0(SUM_AB[5]), .B1(N134), .Y(N438) );
  AOI22X1TF U884 ( .A0(N127), .A1(\INTADD_0_SUM[2] ), .B0(SUM_AB[3]), .B1(N135), .Y(N421) );
  NAND3X1TF U885 ( .A(N905), .B(N219), .C(N218), .Y(N674) );
  NAND4BX1TF U886 ( .AN(N844), .B(N214), .C(N845), .D(N213), .Y(N680) );
  AOI2BB2X1TF U887 ( .B0(N114), .B1(C152_DATA4_2), .A0N(N162), .A1N(N929), .Y(
        N213) );
  OAI2BB1X1TF U888 ( .A0N(N114), .A1N(C152_DATA4_10), .B0(N220), .Y(N672) );
  NAND3X1TF U889 ( .A(N872), .B(N873), .C(N216), .Y(N677) );
  OAI2BB2XLTF U890 ( .B0(OFFSET[0]), .B1(N207), .A0N(Y_IN[2]), .A1N(N81), .Y(
        C2_Z_2) );
  AOI2BB2X1TF U891 ( .B0(N224), .B1(DIVISION_REMA[0]), .A0N(N150), .A1N(N86), 
        .Y(N227) );
  OAI222X1TF U892 ( .A0(N84), .A1(N179), .B0(N86), .B1(N649), .C0(N104), .C1(
        N161), .Y(FOUT[10]) );
  OAI222X1TF U893 ( .A0(N104), .A1(N529), .B0(N86), .B1(N168), .C0(N159), .C1(
        N84), .Y(FOUT[9]) );
  NAND2X1TF U894 ( .A(N152), .B(N170), .Y(N373) );
  NAND3X1TF U895 ( .A(STEP[2]), .B(STEP[3]), .C(N643), .Y(N940) );
  NAND3X1TF U896 ( .A(N546), .B(N385), .C(N635), .Y(N648) );
  NOR4XLTF U897 ( .A(N763), .B(N618), .C(N802), .D(N648), .Y(N266) );
  AOI222XLTF U898 ( .A0(STEP[2]), .A1(N153), .B0(N121), .B1(N170), .C0(N151), 
        .C1(N122), .Y(N264) );
  NAND3X1TF U899 ( .A(N266), .B(N364), .C(N634), .Y(N620) );
  NAND2X1TF U900 ( .A(Y_IN[1]), .B(Y_IN[0]), .Y(N318) );
  AOI2BB1X1TF U901 ( .A0N(N106), .A1N(N273), .B0(Y_IN[4]), .Y(N271) );
  AOI2BB1X1TF U902 ( .A0N(X_IN[7]), .A1N(N277), .B0(Y_IN[6]), .Y(N275) );
  NAND2X1TF U903 ( .A(MODE_TYPE[0]), .B(N315), .Y(N764) );
  AO22X1TF U904 ( .A0(X_IN[4]), .A1(N738), .B0(N93), .B1(N318), .Y(N288) );
  NAND2X1TF U905 ( .A(N105), .B(N731), .Y(N290) );
  AOI2BB1X1TF U906 ( .A0N(N294), .A1N(X_IN[6]), .B0(Y_IN[4]), .Y(N292) );
  AOI2BB1X1TF U907 ( .A0N(N298), .A1N(X_IN[8]), .B0(Y_IN[6]), .Y(N296) );
  NAND2X1TF U908 ( .A(N163), .B(N186), .Y(N617) );
  NAND4BX1TF U909 ( .AN(N381), .B(N316), .C(N804), .D(N364), .Y(N725) );
  NAND2X1TF U910 ( .A(N839), .B(N162), .Y(N847) );
  NAND2X1TF U911 ( .A(N858), .B(N181), .Y(N867) );
  NOR2BX1TF U912 ( .AN(N892), .B(OPER_B[7]), .Y(N895) );
  NAND2X1TF U913 ( .A(N895), .B(N165), .Y(N908) );
  NAND2X1TF U914 ( .A(N923), .B(N166), .Y(N936) );
  NAND2X1TF U915 ( .A(N343), .B(N180), .Y(N348) );
  NAND2X1TF U916 ( .A(N907), .B(N74), .Y(N958) );
  NAND2X1TF U917 ( .A(N566), .B(N958), .Y(N939) );
  NAND2X1TF U918 ( .A(N967), .B(N379), .Y(N574) );
  NAND3X1TF U919 ( .A(N92), .B(N91), .C(N90), .Y(N592) );
  NOR2BX1TF U920 ( .AN(N574), .B(N606), .Y(N571) );
  NAND2X1TF U921 ( .A(PRE_WORK), .B(N354), .Y(N953) );
  NAND2X1TF U922 ( .A(N606), .B(N824), .Y(N347) );
  NAND2X1TF U923 ( .A(N223), .B(N959), .Y(N366) );
  NAND3X1TF U924 ( .A(SIGN_Y), .B(N74), .C(N906), .Y(N825) );
  NAND2X1TF U925 ( .A(N862), .B(N855), .Y(N868) );
  NAND2X1TF U926 ( .A(N881), .B(N882), .Y(N893) );
  NAND2X1TF U927 ( .A(N897), .B(N898), .Y(N909) );
  NAND2X1TF U928 ( .A(N915), .B(N917), .Y(N933) );
  NAND3X1TF U929 ( .A(N606), .B(N603), .C(N167), .Y(N601) );
  NAND2X1TF U930 ( .A(N414), .B(N413), .Y(N422) );
  NAND2X1TF U931 ( .A(N433), .B(N432), .Y(N443) );
  NAND2X1TF U932 ( .A(N453), .B(N452), .Y(N462) );
  NAND2X1TF U933 ( .A(N499), .B(N498), .Y(N1014) );
  AOI222XLTF U934 ( .A0(XTEMP[11]), .A1(N139), .B0(XTEMP[11]), .B1(N497), .C0(
        N139), .C1(N497), .Y(N355) );
  XOR2X1TF U935 ( .A(X_IN[12]), .B(N355), .Y(N360) );
  NAND3X1TF U936 ( .A(N567), .B(POST_WORK), .C(N603), .Y(N376) );
  NAND3BX1TF U937 ( .AN(N366), .B(N949), .C(N967), .Y(N599) );
  NAND3X1TF U938 ( .A(N610), .B(N367), .C(N599), .Y(N943) );
  NAND2X1TF U939 ( .A(N119), .B(N393), .Y(N380) );
  NAND3X1TF U940 ( .A(N383), .B(N122), .C(DP_OP_333_124_4748_N57), .Y(N639) );
  NOR2BX1TF U941 ( .AN(N635), .B(N944), .Y(N543) );
  NAND2X1TF U942 ( .A(N800), .B(SUM_AB[8]), .Y(N424) );
  NAND4X1TF U943 ( .A(N427), .B(N426), .C(N425), .D(N424), .Y(N428) );
  NAND4X1TF U944 ( .A(N438), .B(N437), .C(N436), .D(N435), .Y(N439) );
  NAND4X1TF U945 ( .A(N448), .B(N447), .C(N446), .D(N445), .Y(N449) );
  OAI2BB1X1TF U946 ( .A0N(DIVISION_HEAD[10]), .A1N(N471), .B0(N451), .Y(N713)
         );
  AOI2BB2X1TF U947 ( .B0(X_IN[9]), .B1(N478), .A0N(N478), .A1N(X_IN[9]), .Y(
        N483) );
  NAND3X1TF U948 ( .A(N126), .B(N529), .C(N483), .Y(N479) );
  AOI2BB1X1TF U949 ( .A0N(N509), .A1N(N483), .B0(N513), .Y(N484) );
  AOI2BB2X1TF U950 ( .B0(N487), .B1(N502), .A0N(N502), .A1N(N487), .Y(N494) );
  AOI2BB1X1TF U951 ( .A0N(N509), .A1N(N494), .B0(N513), .Y(N495) );
  AOI2BB2X1TF U952 ( .B0(N139), .B1(N497), .A0N(N497), .A1N(N139), .Y(N510) );
  OAI2BB2XLTF U953 ( .B0(N502), .B1(N609), .A0N(XTEMP[12]), .A1N(N95), .Y(N503) );
  AOI2BB1X1TF U954 ( .A0N(N509), .A1N(N510), .B0(N513), .Y(N511) );
  AOI2BB1X1TF U955 ( .A0N(DIVISION_REMA[2]), .A1N(N518), .B0(DIVISION_HEAD[6]), 
        .Y(N516) );
  OA21XLTF U956 ( .A0(N155), .A1(DIVISION_REMA[4]), .B0(N520), .Y(N522) );
  OA21XLTF U957 ( .A0(N160), .A1(DIVISION_REMA[6]), .B0(N524), .Y(N526) );
  OA21XLTF U958 ( .A0(XTEMP[12]), .A1(N536), .B0(N649), .Y(N535) );
  NAND4X1TF U959 ( .A(N546), .B(N545), .C(N639), .D(N544), .Y(N557) );
  NAND3X1TF U960 ( .A(N552), .B(N551), .C(N550), .Y(N553) );
  NAND3X1TF U961 ( .A(N757), .B(N560), .C(N559), .Y(N561) );
  NAND3X1TF U962 ( .A(N567), .B(N603), .C(N823), .Y(N573) );
  NAND4X1TF U963 ( .A(N569), .B(N568), .C(N640), .D(N573), .Y(N570) );
  NAND2X1TF U964 ( .A(N185), .B(N164), .Y(N591) );
  NOR4XLTF U965 ( .A(\RSHT_BITS[3] ), .B(N90), .C(N615), .D(N591), .Y(N572) );
  NAND2X1TF U966 ( .A(N580), .B(N590), .Y(N587) );
  NAND2X1TF U967 ( .A(N92), .B(N91), .Y(N589) );
  AOI2BB2X1TF U968 ( .B0(N597), .B1(N164), .A0N(N591), .A1N(N593), .Y(N585) );
  NAND4X1TF U969 ( .A(N98), .B(N635), .C(N634), .D(N633), .Y(N636) );
  NAND4X1TF U970 ( .A(N641), .B(N640), .C(N639), .D(N644), .Y(N697) );
  NAND3X1TF U971 ( .A(N757), .B(N653), .C(N652), .Y(N654) );
  AO22X1TF U972 ( .A0(DIVISION_REMA[4]), .A1(N736), .B0(N197), .B1(N791), .Y(
        N744) );
  AOI2BB1X1TF U973 ( .A0N(X_IN[1]), .A1N(N765), .B0(N764), .Y(N768) );
  NAND4X1TF U974 ( .A(N795), .B(N794), .C(N793), .D(N792), .Y(N796) );
  OAI221XLTF U975 ( .A0(\INDEX[2] ), .A1(N90), .B0(N124), .B1(\RSHT_BITS[3] ), 
        .C0(N818), .Y(N819) );
  OAI221XLTF U976 ( .A0(N129), .A1(N185), .B0(N163), .B1(N92), .C0(N820), .Y(
        N836) );
  NAND2X1TF U977 ( .A(N904), .B(N876), .Y(N871) );
  NAND2BX1TF U978 ( .AN(N821), .B(N871), .Y(N891) );
  NAND2X1TF U979 ( .A(N835), .B(N967), .Y(N877) );
  NAND3X1TF U980 ( .A(SIGN_Y), .B(N74), .C(N225), .Y(N843) );
  OAI2BB1X1TF U981 ( .A0N(N960), .A1N(N836), .B0(N835), .Y(N920) );
  NAND3X1TF U982 ( .A(N74), .B(N182), .C(N61), .Y(N975) );
  NAND4X1TF U983 ( .A(N225), .B(N182), .C(N61), .D(N965), .Y(N845) );
  NAND2X1TF U984 ( .A(N904), .B(N920), .Y(N938) );
  NAND2X1TF U985 ( .A(N941), .B(N946), .Y(N947) );
  NAND2X1TF U986 ( .A(N979), .B(N978), .Y(N668) );
  NAND2X1TF U987 ( .A(N982), .B(N981), .Y(N667) );
  NAND2X1TF U988 ( .A(SUM_AB[3]), .B(N88), .Y(N983) );
  NAND2X1TF U989 ( .A(N988), .B(N987), .Y(N665) );
  NAND2X1TF U990 ( .A(SUM_AB[5]), .B(N88), .Y(N989) );
  NAND2X1TF U991 ( .A(N994), .B(N993), .Y(N663) );
  NAND2X1TF U992 ( .A(SUM_AB[7]), .B(N88), .Y(N995) );
  NAND2X1TF U993 ( .A(N1000), .B(N999), .Y(N661) );
  NAND2X1TF U994 ( .A(SUM_AB[9]), .B(N88), .Y(N1001) );
  NAND2X1TF U995 ( .A(N1006), .B(N1005), .Y(N659) );
  NAND2X1TF U996 ( .A(SUM_AB[11]), .B(N88), .Y(N1007) );
endmodule


module SERIAL_CPU_8BIT_VG ( CLK, ENABLE, RST_N, START, I_DATAIN, D_DATAIN, 
        CPU_WAIT, IS_I_ADDR, NXT, I_ADDR, D_ADDR, D_WE, D_DATAOUT, IO_STATUS, 
        IO_DATAINA, IO_DATAINB, IO_DATAOUTA, IO_DATAOUTB, IO_OFFSET, I_PC, 
        I_REG_C, \IO_CONTROL[15] , \IO_CONTROL[14] , \IO_CONTROL[13] , 
        \IO_CONTROL[12] , \IO_CONTROL[11] , \IO_CONTROL[10] , \IO_CONTROL[9] , 
        \IO_CONTROL[8] , \IO_CONTROL[7] , \IO_CONTROL[6] , \IO_CONTROL[5]_BAR , 
        \IO_CONTROL[4] , \IO_CONTROL[3] , \IO_CONTROL[2] , \IO_CONTROL[1] , 
        \IO_CONTROL[0]  );
  input [7:0] I_DATAIN;
  input [7:0] D_DATAIN;
  output [1:0] NXT;
  output [9:0] I_ADDR;
  output [9:0] D_ADDR;
  output [7:0] D_DATAOUT;
  input [15:0] IO_STATUS;
  input [15:0] IO_DATAINA;
  input [15:0] IO_DATAINB;
  output [15:0] IO_DATAOUTA;
  output [15:0] IO_DATAOUTB;
  output [15:0] IO_OFFSET;
  output [5:0] I_PC;
  output [5:0] I_REG_C;
  input CLK, ENABLE, RST_N, START, CPU_WAIT;
  output IS_I_ADDR, D_WE, \IO_CONTROL[15] , \IO_CONTROL[14] , \IO_CONTROL[13] ,
         \IO_CONTROL[12] , \IO_CONTROL[11] , \IO_CONTROL[10] , \IO_CONTROL[9] ,
         \IO_CONTROL[8] , \IO_CONTROL[7] , \IO_CONTROL[6] ,
         \IO_CONTROL[5]_BAR , \IO_CONTROL[4] , \IO_CONTROL[3] ,
         \IO_CONTROL[2] , \IO_CONTROL[1] , \IO_CONTROL[0] ;
  wire   N89, N90, N91, N92, N93, N94, N95, N96, N97, N1356, N1357, N1358,
         N1359, N1360, N1361, N1362, N1363, \IO_CONTROL[5] , N1364, N1365,
         N1366, N1367, N1368, N1369, N1370, N1371, N1372, N1373, N1374, N1375,
         \GR[7][15] , \GR[7][14] , \GR[7][13] , \GR[7][12] , \GR[7][11] ,
         \GR[7][10] , \GR[7][9] , \GR[7][8] , \GR[7][7] , \GR[7][6] ,
         \GR[7][5] , \GR[7][4] , \GR[7][3] , \GR[7][2] , \GR[7][1] ,
         \GR[7][0] , \GR[6][15] , \GR[6][14] , \GR[6][13] , \GR[6][12] ,
         \GR[6][11] , \GR[6][10] , \GR[6][9] , \GR[6][8] , \GR[6][7] ,
         \GR[6][6] , \GR[6][5] , \GR[6][4] , \GR[6][3] , \GR[6][2] ,
         \GR[6][1] , \GR[6][0] , \GR[5][15] , \GR[5][14] , \GR[5][13] ,
         \GR[5][12] , \GR[5][11] , \GR[5][10] , \GR[5][9] , \GR[5][8] ,
         \GR[5][7] , \GR[5][6] , \GR[5][5] , \GR[5][4] , \GR[5][3] ,
         \GR[5][2] , \GR[5][1] , \GR[5][0] , \GR[0][15] , \GR[0][14] ,
         \GR[0][13] , \GR[0][12] , \GR[0][11] , \GR[0][10] , \GR[0][9] ,
         \GR[0][8] , \GR[0][7] , \GR[0][6] , \GR[0][5] , \GR[0][4] ,
         \GR[0][3] , \GR[0][2] , \GR[0][1] , \GR[0][0] , N157, N158, N159,
         N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172,
         N173, N174, N175, N176, N177, N199, N200, N201, N202, N203, N204,
         N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N239,
         N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250,
         N251, N252, N253, N254, CF_BUF, N449, N450, N451, N452, N453, N454,
         N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, N465,
         N483, N484, N485, N486, N487, N488, N489, N490, N491, N492, N493,
         N494, N495, N496, N497, N498, N499, N567, N568, ZF, NF, CF, N595,
         N259, N260, N279, N424, N426, N428, N430, N432, N434, N436, N438,
         N440, N442, N444, N446, N448, N4500, N4520, N4540, N4550, N4560,
         N4570, N4590, N4600, N4610, N4620, N4630, N4640, N4650, N466, N467,
         N468, N469, N470, N471, N472, N473, N474, N475, N476, N477, N478,
         N479, N480, N481, N482, N4830, N4840, N4850, N4860, N4870, N4880,
         N4890, N4900, N4910, N4920, N4930, N4940, N4950, N4960, N4970, N4980,
         N4990, N500, N501, N502, N503, N504, N505, N506, N507, N508, N509,
         N510, N511, N512, N513, N514, N517, N518, N519, N520, N522, N523,
         N524, N526, N552, N5670, N572, N573, N574, N575, N577, N578, N579,
         N580, N581, N582, N583, N606, N717, N721, N722, N724, N725, N726,
         N776, N777, N832, N833, N834, N835, N836, N837, N838, N839, N840,
         N841, N842, N843, N844, N845, N846, N847, N848, N849, N850, N851,
         N852, N853, N854, N855, N856, N857, N858, N859, N860, N861, N862,
         N863, N864, N865, N866, N867, N868, N869, N870, N871, N872, N873,
         N874, N875, N876, N877, N878, N879, N880, N881, N882, N883, N884,
         N885, N886, N887, N888, N889, N890, N891, N892, N893, N894, N895,
         N896, N897, N898, N899, N900, N901, N902, N903, N904, N905, N906,
         N907, N908, N909, N910, N911, N912, N913, N914, N915, N916, N917,
         N918, N919, N920, N921, N922, N923, N924, N925, N926, N927, N928,
         N929, N930, N931, N932, N933, N934, N935, N936, N937, N938, N939,
         N940, N941, N942, N943, N944, N945, N946, N947, N948, N949, N950,
         N951, N952, N953, N954, N955, N956, N957, N958, N959, N960, N961,
         N962, ADD_X_300_3_N22, ADD_X_300_3_N21, ADD_X_300_3_N20,
         ADD_X_300_3_N19, ADD_X_300_3_N18, ADD_X_300_3_N17, ADD_X_300_3_N16,
         ADD_X_300_3_N15, ADD_X_300_3_N14, ADD_X_300_3_N13, ADD_X_300_3_N12,
         ADD_X_300_3_N11, ADD_X_300_3_N10, ADD_X_300_3_N9, ADD_X_300_3_N8,
         ADD_X_300_3_N7, ADD_X_300_3_N6, ADD_X_300_3_N5, ADD_X_300_3_N4,
         ADD_X_300_3_N3, ADD_X_300_3_N2, SUB_X_300_4_N16, SUB_X_300_4_N15,
         SUB_X_300_4_N14, SUB_X_300_4_N13, SUB_X_300_4_N12, SUB_X_300_4_N11,
         SUB_X_300_4_N10, SUB_X_300_4_N9, SUB_X_300_4_N8, SUB_X_300_4_N7,
         SUB_X_300_4_N6, SUB_X_300_4_N5, SUB_X_300_4_N4, SUB_X_300_4_N3,
         SUB_X_300_4_N2, SUB_X_300_4_N1, N1, N2, N3, N4, N5, N6, N7, N8, N9,
         N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23,
         N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, N189, N191, N193, N195, N197, N198,
         N1990, N2000, N2010, N2030, N2050, N2070, N2090, N2100, N2110, N2120,
         N2130, N2140, N216, N217, N218, N220, N221, N222, N223, N224, N225,
         N226, N227, N228, N229, N230, N231, N232, N233, N234, N235, N236,
         N237, N238, N2390, N2400, N2410, N2420, N2430, N2440, N2450, N2460,
         N2470, N2480, N2490, N2500, N2510, N2520, N2530, N2540, N255, N256,
         N257, N258, N261, N262, N263, N264, N265, N266, N267, N268, N269,
         N270, N271, N272, N273, N274, N275, N276, N277, N278, N280, N281,
         N282, N283, N284, N285, N286, N288, N290, N292, N293, N294, N295,
         N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, N306,
         N307, N308, N309, N310, N311, N332, N333, N334, N335, N336, N337,
         N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, N348,
         N349, N350, N351, N352, N353, N354, N355, N356, N357, N358, N359,
         N360, N361, N362, N363, N364, N365, N366, N367, N368, N369, N370,
         N371, N372, N373, N374, N375, N376, N377, N378, N379, N380, N381,
         N382, N383, N384, N385, N386, N387, N388, N389, N390, N391, N392,
         N393, N394, N395, N396, N397, N398, N399, N400, N401, N402, N403,
         N404, N405, N406, N407, N408, N409, N410, N411, N412, N413, N414,
         N415, N416, N417, N418, N419, N420, N421, N422, N423, N425, N427,
         N429, N431, N433, N435, N437, N439, N441, N443, N445, N447, N4490,
         N4510, N4530, N4580, N516, N521, N525, N527, N528, N529, N530, N531,
         N532, N533, N534, N535, N536, N537, N538, N539, N540, N541, N542,
         N543, N544, N545, N546, N547, N548, N549, N550, N551, N553, N554,
         N555, N556, N557, N558, N559, N560, N561, N562, N563, N564, N565,
         N566, N5680, N569, N570, N571, N576, N584, N585, N586, N587, N588,
         N589, N590, N591, N592, N593, N594, N5950, N596, N597, N598, N599,
         N600, N601, N602, N603, N604, N605, N607, N608, N609, N610, N611,
         N612, N613, N614, N615, N616, N617, N618, N619, N620, N621, N622,
         N623, N624, N625, N626, N627, N628, N629, N630, N631, N632, N633,
         N634, N635, N636, N637, N638, N639, N640, N641, N642, N643, N644,
         N645, N646, N647, N648, N649, N650, N651, N652, N653, N654, N655,
         N656, N657, N658, N659, N660, N661, N662, N663, N664, N665, N666,
         N667, N668, N669, N670, N671, N672, N673, N674, N675, N676, N677,
         N678, N679, N680, N681, N682, N683, N684, N685, N686, N687, N688,
         N689, N690, N691, N692, N693, N694, N695, N696, N697, N698, N699,
         N700, N701, N702, N703, N704, N705, N706, N707, N708, N709, N710,
         N711, N712, N713, N714, N715, N716, N718, N719, N720, N723, N727,
         N728, N729, N730, N731, N732, N733, N734, N735, N736, N737, N738,
         N739, N740, N741, N742, N743, N744, N745, N746, N747, N748, N749,
         N750, N751, N752, N753, N754, N755, N756, N757, N758, N759, N760,
         N761, N762, N763, N764, N765, N766, N767, N768, N769, N770, N771,
         N772, N773, N774, N775, N778, N779, N780, N781, N782, N783, N784,
         N785, N786, N787, N788, N789, N790, N791, N792, N793, N794, N795,
         N796, N797, N798, N799, N800, N801, N802, N803, N804, N805, N806,
         N807, N808, N809, N810, N811, N812, N813, N814, N815, N816, N817,
         N818, N819, N820, N821, N822, N823, N824, N825, N826, N827, N828,
         N829, N830, N831, N963, N964, N965, N966, N967, N968, N969, N970,
         N971, N972, N973, N974, N975, N976, N977, N978, N979, N980, N981,
         N982, N983, N984, N985, N986, N987, N988, N989, N990, N991, N992,
         N993, N994, N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003,
         N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013,
         N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023,
         N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1031, N1032, N1033,
         N1034, N1035, N1036, N1037, N1038, N1039, N1040, N1041, N1042, N1043,
         N1044, N1045, N1046, N1047, N1048, N1049, N1050, N1051, N1052, N1053,
         N1054, N1055, N1056, N1057, N1058, N1059, N1060, N1061, N1062, N1063,
         N1064, N1065, N1066, N1067, N1068, N1069, N1070, N1071, N1072, N1073,
         N1074, N1075, N1076, N1077, N1078, N1079, N1080, N1081, N1082, N1083,
         N1084, N1085, N1086, N1087, N1088, N1089, N1090, N1091, N1092, N1093,
         N1094, N1095, N1096, N1097, N1098, N1099, N1100, N1101, N1102, N1103,
         N1104, N1105, N1106, N1107, N1108, N1109, N1110, N1111, N1112, N1113,
         N1114, N1115, N1116, N1117, N1118, N1119, N1120, N1121, N1122, N1123,
         N1124, N1125, N1126, N1127, N1128, N1129, N1130, N1131, N1132, N1133,
         N1134, N1135, N1136, N1137, N1138, N1139, N1140, N1141, N1142, N1143,
         N1144, N1145, N1146, N1147, N1148, N1149, N1150, N1151, N1152, N1153,
         N1154, N1155, N1156, N1157, N1158, N1159, N1160, N1161, N1162, N1163,
         N1164, N1165, N1166, N1167, N1168, N1169, N1170, N1171, N1172, N1173,
         N1174, N1175, N1176, N1177, N1178, N1179, N1180, N1181, N1182, N1183,
         N1184, N1185, N1186, N1187, N1188, N1189, N1190, N1191, N1192, N1193,
         N1194, N1195, N1196, N1197, N1198, N1199, N1200, N1201, N1202, N1203,
         N1204, N1205, N1206, N1207, N1208, N1209, N1210, N1211, N1212, N1213,
         N1214, N1215, N1216, N1217, N1218, N1219, N1220, N1221, N1222, N1223,
         N1224, N1225, N1226, N1227, N1228, N1229, N1230, N1231, N1232, N1233,
         N1234, N1235, N1236, N1237, N1238, N1239, N1240, N1241, N1242, N1243,
         N1244, N1245, N1246, N1247, N1248, N1249, N1250, N1251, N1252, N1253,
         N1254, N1255, N1256, N1257, N1258, N1259, N1260, N1261, N1262, N1263,
         N1264, N1265, N1266, N1267, N1268, N1269, N1270, N1271, N1272, N1273,
         N1274, N1275, N1276, N1277, N1278, N1279, N1280, N1281, N1282, N1283,
         N1284, N1285, N1286, N1287, N1288, N1289, N1290, N1291, N1292, N1293,
         N1294, N1295, N1296, N1297, N1298, N1299, N1300, N1301, N1302, N1303,
         N1304, N1305, N1306, N1307, N1308, N1309, N1310, N1311, N1312, N1313,
         N1314, N1315, N1316, N1317, N1318, N1319, N1320, N1321, N1322, N1323,
         N1324, N1325, N1326, N1327, N1328, N1329, N1330, N1331, N1332, N1333,
         N1334, N1335, N1336, N1337, N1338, N1339, N1340, N1341, N1342, N1343,
         N1344, N1345, N1346, N1347, N1348, N1349, N1350, N1351, N1352, N1353,
         N1354, N1355;
  wire   [15:9] REG_C;
  wire   [3:1] CODE_TYPE;
  wire   [3:1] STATE;
  wire   [3:0] NEXT_STATE;
  wire   [15:0] REG_A;
  wire   [15:0] REG_B;
  wire   [15:0] SMDR;

  CLKINVX6TF U412 ( .A(RST_N), .Y(N606) );
  AFCSIHCONX2TF \add_x_300_3/U17  ( .A(REG_A[2]), .B(REG_B[2]), .CS(
        ADD_X_300_3_N21), .S(N451), .CO0N(ADD_X_300_3_N20), .CO1N(
        ADD_X_300_3_N19) );
  AFCSHCINX2TF \add_x_300_3/U16  ( .CI1N(ADD_X_300_3_N19), .B(REG_A[3]), .A(
        REG_B[3]), .CI0N(ADD_X_300_3_N20), .CS(ADD_X_300_3_N21), .CO1(
        ADD_X_300_3_N17), .CO0(ADD_X_300_3_N18), .S(N452) );
  AFCSIHCONX2TF \add_x_300_3/U14  ( .A(REG_A[4]), .B(REG_B[4]), .CS(
        ADD_X_300_3_N16), .S(N453), .CO0N(ADD_X_300_3_N15), .CO1N(
        ADD_X_300_3_N14) );
  AFCSHCINX2TF \add_x_300_3/U13  ( .CI1N(ADD_X_300_3_N14), .B(REG_A[5]), .A(
        REG_B[5]), .CI0N(ADD_X_300_3_N15), .CS(ADD_X_300_3_N16), .CO1(
        ADD_X_300_3_N12), .CO0(ADD_X_300_3_N13), .S(N454) );
  CMPR32X2TF \add_x_300_3/U11  ( .A(REG_A[6]), .B(REG_B[6]), .C(
        ADD_X_300_3_N11), .CO(ADD_X_300_3_N10), .S(N455) );
  CMPR32X2TF \add_x_300_3/U10  ( .A(REG_A[7]), .B(REG_B[7]), .C(
        ADD_X_300_3_N10), .CO(ADD_X_300_3_N9), .S(N456) );
  CMPR32X2TF \add_x_300_3/U9  ( .A(REG_A[8]), .B(REG_B[8]), .C(ADD_X_300_3_N9), 
        .CO(ADD_X_300_3_N8), .S(N457) );
  CMPR32X2TF \add_x_300_3/U8  ( .A(REG_A[9]), .B(REG_B[9]), .C(ADD_X_300_3_N8), 
        .CO(ADD_X_300_3_N7), .S(N458) );
  CMPR32X2TF \add_x_300_3/U7  ( .A(REG_A[10]), .B(REG_B[10]), .C(
        ADD_X_300_3_N7), .CO(ADD_X_300_3_N6), .S(N459) );
  CMPR32X2TF \add_x_300_3/U6  ( .A(REG_A[11]), .B(REG_B[11]), .C(
        ADD_X_300_3_N6), .CO(ADD_X_300_3_N5), .S(N460) );
  CMPR32X2TF \add_x_300_3/U5  ( .A(REG_A[12]), .B(REG_B[12]), .C(
        ADD_X_300_3_N5), .CO(ADD_X_300_3_N4), .S(N461) );
  CMPR32X2TF \add_x_300_3/U4  ( .A(REG_A[13]), .B(REG_B[13]), .C(
        ADD_X_300_3_N4), .CO(ADD_X_300_3_N3), .S(N462) );
  CMPR32X2TF \add_x_300_3/U3  ( .A(REG_A[14]), .B(REG_B[14]), .C(
        ADD_X_300_3_N3), .CO(ADD_X_300_3_N2), .S(N463) );
  DFFRX2TF \state_reg[2]  ( .D(NEXT_STATE[2]), .CK(CLK), .RN(RST_N), .Q(
        STATE[2]), .QN(N348) );
  DFFRX2TF \state_reg[1]  ( .D(NEXT_STATE[1]), .CK(CLK), .RN(RST_N), .Q(
        STATE[1]), .QN(N375) );
  DFFRX2TF \state_reg[0]  ( .D(NEXT_STATE[0]), .CK(CLK), .RN(RST_N), .QN(N552)
         );
  DFFRX2TF \state_reg[3]  ( .D(NEXT_STATE[3]), .CK(CLK), .RN(RST_N), .Q(
        STATE[3]) );
  DFFSX2TF \pc_reg[2]  ( .D(N725), .CK(CLK), .SN(RST_N), .Q(N373), .QN(
        I_ADDR[3]) );
  DFFRX2TF \id_ir_reg[7]  ( .D(N507), .CK(CLK), .RN(RST_N), .Q(N372), .QN(N260) );
  DFFRX2TF \id_ir_reg[4]  ( .D(N510), .CK(CLK), .RN(RST_N), .Q(N92), .QN(N371)
         );
  DFFRX2TF \id_ir_reg[0]  ( .D(N514), .CK(CLK), .RN(RST_N), .Q(N95), .QN(N370)
         );
  DFFRX2TF \id_ir_reg[8]  ( .D(N524), .CK(CLK), .RN(RST_N), .Q(N89), .QN(N369)
         );
  DFFRX2TF zf_reg ( .D(N4570), .CK(CLK), .RN(RST_N), .Q(ZF), .QN(N368) );
  DFFRX2TF nf_reg ( .D(N4560), .CK(CLK), .RN(RST_N), .Q(NF), .QN(N367) );
  DFFSX2TF \pc_reg[7]  ( .D(N717), .CK(CLK), .SN(RST_N), .Q(N366), .QN(
        I_ADDR[8]) );
  DFFSX2TF \pc_reg[5]  ( .D(N722), .CK(CLK), .SN(RST_N), .Q(N365), .QN(
        I_ADDR[6]) );
  DFFSX2TF \pc_reg[3]  ( .D(N724), .CK(CLK), .SN(RST_N), .Q(N364), .QN(
        I_ADDR[4]) );
  DFFRX2TF \reg_B_reg[14]  ( .D(N4600), .CK(CLK), .RN(RST_N), .Q(REG_B[14]), 
        .QN(N573) );
  DFFRX2TF \reg_A_reg[6]  ( .D(N4840), .CK(CLK), .RN(RST_N), .Q(REG_A[6]), 
        .QN(N363) );
  DFFRX2TF \reg_A_reg[4]  ( .D(N4860), .CK(CLK), .RN(RST_N), .Q(REG_A[4]), 
        .QN(N362) );
  DFFRX2TF \reg_A_reg[5]  ( .D(N4850), .CK(CLK), .RN(RST_N), .Q(REG_A[5]), 
        .QN(N361) );
  DFFRX2TF \reg_B_reg[3]  ( .D(N471), .CK(CLK), .RN(RST_N), .Q(REG_B[3]), .QN(
        N360) );
  DFFRX2TF \reg_B_reg[2]  ( .D(N472), .CK(CLK), .RN(RST_N), .Q(REG_B[2]), .QN(
        N356) );
  DFFRX2TF \id_ir_reg[5]  ( .D(N509), .CK(CLK), .RN(RST_N), .Q(N93), .QN(N353)
         );
  DFFRX2TF \id_ir_reg[1]  ( .D(N513), .CK(CLK), .RN(RST_N), .Q(N96), .QN(N352)
         );
  DFFRX2TF \id_ir_reg[9]  ( .D(N523), .CK(CLK), .RN(RST_N), .Q(N90), .QN(N351)
         );
  DFFRX2TF \reg_A_reg[15]  ( .D(N475), .CK(CLK), .RN(RST_N), .Q(REG_A[15]), 
        .QN(N350) );
  DFFRX2TF \reg_A_reg[13]  ( .D(N477), .CK(CLK), .RN(RST_N), .Q(REG_A[13]), 
        .QN(N345) );
  DFFRX2TF \reg_A_reg[10]  ( .D(N480), .CK(CLK), .RN(RST_N), .Q(REG_A[10]), 
        .QN(N344) );
  DFFRX2TF \reg_A_reg[7]  ( .D(N4830), .CK(CLK), .RN(RST_N), .Q(REG_A[7]), 
        .QN(N343) );
  DFFRX2TF \reg_A_reg[3]  ( .D(N4870), .CK(CLK), .RN(RST_N), .Q(REG_A[3]), 
        .QN(N342) );
  DFFRX2TF \reg_A_reg[8]  ( .D(N482), .CK(CLK), .RN(RST_N), .Q(REG_A[8]), .QN(
        N341) );
  DFFRX2TF \reg_A_reg[9]  ( .D(N481), .CK(CLK), .RN(RST_N), .Q(REG_A[9]), .QN(
        N340) );
  DFFRX2TF \reg_A_reg[2]  ( .D(N4880), .CK(CLK), .RN(RST_N), .Q(REG_A[2]), 
        .QN(N339) );
  DFFRX2TF \reg_A_reg[11]  ( .D(N479), .CK(CLK), .RN(RST_N), .Q(REG_A[11]), 
        .QN(N338) );
  DFFRX2TF \id_ir_reg[6]  ( .D(N508), .CK(CLK), .RN(RST_N), .Q(N94), .QN(N337)
         );
  DFFRX2TF \id_ir_reg[2]  ( .D(N512), .CK(CLK), .RN(RST_N), .Q(N97), .QN(N336)
         );
  DFFRX2TF \id_ir_reg[10]  ( .D(N522), .CK(CLK), .RN(RST_N), .Q(N91), .QN(N335) );
  DFFRX2TF \reg_A_reg[14]  ( .D(N476), .CK(CLK), .RN(RST_N), .Q(REG_A[14]), 
        .QN(N334) );
  DFFRX2TF \reg_A_reg[12]  ( .D(N478), .CK(CLK), .RN(RST_N), .Q(REG_A[12]), 
        .QN(N333) );
  DFFRX2TF \reg_A_reg[1]  ( .D(N4890), .CK(CLK), .RN(RST_N), .Q(REG_A[1]), 
        .QN(N332) );
  DFFRX2TF \id_ir_reg[14]  ( .D(N518), .CK(CLK), .RN(RST_N), .Q(CODE_TYPE[3]), 
        .QN(N359) );
  TLATXLTF cf_buf_reg ( .G(N567), .D(N568), .Q(CF_BUF) );
  TLATXLTF \nxt_reg[0]  ( .G(N157), .D(N158), .Q(NXT[0]) );
  TLATXLTF \nxt_reg[1]  ( .G(N157), .D(N159), .Q(NXT[1]) );
  DFFRX2TF \id_ir_reg[3]  ( .D(N511), .CK(CLK), .RN(RST_N), .QN(N259) );
  DFFSX2TF \pc_reg[8]  ( .D(N776), .CK(CLK), .SN(RST_N), .QN(I_ADDR[9]) );
  DFFSX2TF \pc_reg[6]  ( .D(N721), .CK(CLK), .SN(RST_N), .QN(I_ADDR[7]) );
  DFFSX2TF \pc_reg[1]  ( .D(N726), .CK(CLK), .SN(RST_N), .QN(I_ADDR[2]) );
  DFFSX2TF \pc_reg[0]  ( .D(N777), .CK(CLK), .SN(RST_N), .QN(I_ADDR[1]) );
  DFFRX2TF \reg_B_reg[15]  ( .D(N4590), .CK(CLK), .RN(RST_N), .Q(REG_B[15]), 
        .QN(N572) );
  DFFNSRX2TF \reg_C_reg[12]  ( .D(N448), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        REG_C[12]) );
  DFFNSRX2TF \reg_C_reg[11]  ( .D(N446), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        REG_C[11]) );
  DFFNSRX2TF \reg_C_reg[10]  ( .D(N444), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        REG_C[10]) );
  DFFRX2TF \reg_B_reg[10]  ( .D(N4640), .CK(CLK), .RN(RST_N), .Q(REG_B[10]), 
        .QN(N577) );
  DFFRX2TF \reg_B_reg[12]  ( .D(N4620), .CK(CLK), .RN(RST_N), .Q(REG_B[12]), 
        .QN(N575) );
  DFFRX2TF \reg_B_reg[13]  ( .D(N4610), .CK(CLK), .RN(RST_N), .Q(REG_B[13]), 
        .QN(N574) );
  DFFNSRX2TF \reg_C_reg[15]  ( .D(N4540), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        REG_C[15]) );
  DFFNSRX2TF \reg_C_reg[6]  ( .D(N436), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[7]) );
  DFFNSRX2TF \reg_C_reg[7]  ( .D(N438), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[8]) );
  DFFRX2TF \reg_B_reg[6]  ( .D(N468), .CK(CLK), .RN(RST_N), .Q(REG_B[6]), .QN(
        N581) );
  DFFRX2TF \reg_B_reg[7]  ( .D(N467), .CK(CLK), .RN(RST_N), .Q(REG_B[7]), .QN(
        N580) );
  DFFRX2TF \reg_B_reg[8]  ( .D(N466), .CK(CLK), .RN(RST_N), .Q(REG_B[8]), .QN(
        N579) );
  DFFRX2TF \reg_B_reg[9]  ( .D(N4650), .CK(CLK), .RN(RST_N), .Q(REG_B[9]), 
        .QN(N578) );
  DFFRX2TF \reg_B_reg[5]  ( .D(N469), .CK(CLK), .RN(RST_N), .Q(REG_B[5]), .QN(
        N582) );
  DFFRX2TF \reg_B_reg[4]  ( .D(N470), .CK(CLK), .RN(RST_N), .Q(REG_B[4]), .QN(
        N583) );
  DFFNSRX2TF \reg_C_reg[1]  ( .D(N426), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[2]) );
  DFFNSRX2TF \reg_C_reg[5]  ( .D(N434), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[6]) );
  DFFNSRX2TF \reg_C_reg[4]  ( .D(N432), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[5]) );
  DFFNSRX2TF \reg_C_reg[0]  ( .D(N424), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[1]) );
  DFFNSRX2TF \reg_C_reg[3]  ( .D(N430), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[4]) );
  DFFRX2TF \id_ir_reg[12]  ( .D(N520), .CK(CLK), .RN(RST_N), .Q(CODE_TYPE[1]), 
        .QN(N306) );
  CMPR32X2TF \add_x_300_3/U2  ( .A(REG_A[15]), .B(REG_B[15]), .C(
        ADD_X_300_3_N2), .CO(N465), .S(N464) );
  CMPR32X2TF \add_x_300_3/U18  ( .A(REG_B[1]), .B(REG_A[1]), .C(
        ADD_X_300_3_N22), .CO(ADD_X_300_3_N21), .S(N450) );
  CLKMX2X2TF \add_x_300_3/U12  ( .A(ADD_X_300_3_N13), .B(ADD_X_300_3_N12), 
        .S0(ADD_X_300_3_N16), .Y(ADD_X_300_3_N11) );
  CLKMX2X4TF \add_x_300_3/U15  ( .A(ADD_X_300_3_N18), .B(ADD_X_300_3_N17), 
        .S0(ADD_X_300_3_N21), .Y(ADD_X_300_3_N16) );
  DFFNSRX2TF \reg_C_reg[2]  ( .D(N428), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[3]) );
  CMPR32X2TF \sub_x_300_4/U11  ( .A(N581), .B(REG_A[6]), .C(SUB_X_300_4_N11), 
        .CO(SUB_X_300_4_N10), .S(N489) );
  CMPR32X2TF \sub_x_300_4/U12  ( .A(N582), .B(REG_A[5]), .C(SUB_X_300_4_N12), 
        .CO(SUB_X_300_4_N11), .S(N488) );
  CMPR32X2TF \sub_x_300_4/U6  ( .A(N311), .B(REG_A[11]), .C(SUB_X_300_4_N6), 
        .CO(SUB_X_300_4_N5), .S(N494) );
  ADDFHX1TF \sub_x_300_4/U8  ( .A(N578), .B(REG_A[9]), .CI(SUB_X_300_4_N8), 
        .CO(SUB_X_300_4_N7), .S(N492) );
  CMPR32X2TF \sub_x_300_4/U10  ( .A(N580), .B(REG_A[7]), .C(SUB_X_300_4_N10), 
        .CO(SUB_X_300_4_N9), .S(N490) );
  CMPR32X2TF \sub_x_300_4/U13  ( .A(N583), .B(REG_A[4]), .C(SUB_X_300_4_N13), 
        .CO(SUB_X_300_4_N12), .S(N487) );
  CMPR32X2TF \sub_x_300_4/U14  ( .A(N360), .B(REG_A[3]), .C(SUB_X_300_4_N14), 
        .CO(SUB_X_300_4_N13), .S(N486) );
  CMPR32X2TF \sub_x_300_4/U9  ( .A(N579), .B(REG_A[8]), .C(SUB_X_300_4_N9), 
        .CO(SUB_X_300_4_N8), .S(N491) );
  CMPR32X2TF \sub_x_300_4/U3  ( .A(N573), .B(REG_A[14]), .C(SUB_X_300_4_N3), 
        .CO(SUB_X_300_4_N2), .S(N497) );
  CMPR32X2TF \sub_x_300_4/U15  ( .A(N356), .B(REG_A[2]), .C(SUB_X_300_4_N15), 
        .CO(SUB_X_300_4_N14), .S(N485) );
  CMPR32X2TF \sub_x_300_4/U7  ( .A(N577), .B(REG_A[10]), .C(SUB_X_300_4_N7), 
        .CO(SUB_X_300_4_N6), .S(N493) );
  CMPR32X2TF \sub_x_300_4/U5  ( .A(N575), .B(REG_A[12]), .C(SUB_X_300_4_N5), 
        .CO(SUB_X_300_4_N4), .S(N495) );
  CMPR32X2TF \sub_x_300_4/U4  ( .A(N574), .B(REG_A[13]), .C(SUB_X_300_4_N4), 
        .CO(SUB_X_300_4_N3), .S(N496) );
  DFFNSRXLTF \reg_C_reg[9]  ( .D(N442), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        REG_C[9]) );
  DFFNSRXLTF \reg_C_reg[13]  ( .D(N4500), .CKN(CLK), .SN(1'b1), .RN(1'b1), 
        .QN(N279) );
  DFFNSRXLTF is_i_addr_reg ( .D(N961), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        IS_I_ADDR), .QN(N526) );
  DFFNSRXLTF \reg_C_reg[14]  ( .D(N4520), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        REG_C[14]), .QN(N374) );
  DFFNSRXLTF dw_reg ( .D(N595), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(D_WE) );
  DFFRX2TF \reg_A_reg[0]  ( .D(N4900), .CK(CLK), .RN(RST_N), .Q(REG_A[0]), 
        .QN(N349) );
  DFFSX4TF \id_ir_reg[11]  ( .D(N31), .CK(CLK), .SN(RST_N), .Q(N5670), .QN(
        N634) );
  DFFRX1TF \smdr_reg[7]  ( .D(N4990), .CK(CLK), .RN(RST_N), .Q(SMDR[7]) );
  DFFRX1TF \smdr_reg[0]  ( .D(N506), .CK(CLK), .RN(RST_N), .Q(SMDR[0]) );
  DFFRX1TF \smdr_reg[14]  ( .D(N4920), .CK(CLK), .RN(RST_N), .Q(SMDR[14]) );
  DFFRX1TF \smdr_reg[8]  ( .D(N4980), .CK(CLK), .RN(RST_N), .Q(SMDR[8]) );
  DFFRX1TF \smdr_reg[1]  ( .D(N505), .CK(CLK), .RN(RST_N), .Q(SMDR[1]) );
  DFFRX1TF \smdr_reg[15]  ( .D(N4910), .CK(CLK), .RN(RST_N), .Q(SMDR[15]) );
  DFFRX1TF \smdr_reg[13]  ( .D(N4930), .CK(CLK), .RN(RST_N), .Q(SMDR[13]) );
  DFFRX1TF \smdr_reg[10]  ( .D(N4960), .CK(CLK), .RN(RST_N), .Q(SMDR[10]) );
  DFFRX1TF \smdr_reg[11]  ( .D(N4950), .CK(CLK), .RN(RST_N), .Q(SMDR[11]) );
  DFFRX1TF \smdr_reg[12]  ( .D(N4940), .CK(CLK), .RN(RST_N), .Q(SMDR[12]) );
  DFFRX1TF \smdr_reg[9]  ( .D(N4970), .CK(CLK), .RN(RST_N), .Q(SMDR[9]) );
  DFFRX1TF \smdr_reg[6]  ( .D(N500), .CK(CLK), .RN(RST_N), .Q(SMDR[6]) );
  DFFRX1TF \smdr_reg[5]  ( .D(N501), .CK(CLK), .RN(RST_N), .Q(SMDR[5]) );
  DFFRX1TF \smdr_reg[4]  ( .D(N502), .CK(CLK), .RN(RST_N), .Q(SMDR[4]) );
  DFFRX1TF \smdr_reg[3]  ( .D(N503), .CK(CLK), .RN(RST_N), .Q(SMDR[3]) );
  DFFRX1TF \smdr_reg[2]  ( .D(N504), .CK(CLK), .RN(RST_N), .Q(SMDR[2]) );
  DFFRX1TF cf_reg ( .D(N4550), .CK(CLK), .RN(RST_N), .Q(CF) );
  DFFRX1TF \reg_B_reg[11]  ( .D(N4630), .CK(CLK), .RN(RST_N), .Q(REG_B[11]), 
        .QN(N311) );
  DFFRX1TF \pc_reg[4]  ( .D(N832), .CK(CLK), .RN(RST_N), .Q(I_ADDR[5]) );
  DFFRX1TF \gr_reg[7][13]  ( .D(N835), .CK(CLK), .RN(RST_N), .Q(\GR[7][13] )
         );
  DFFRX1TF \gr_reg[6][13]  ( .D(N843), .CK(CLK), .RN(RST_N), .Q(\GR[6][13] )
         );
  DFFRX1TF \gr_reg[5][13]  ( .D(N851), .CK(CLK), .RN(RST_N), .Q(\GR[5][13] )
         );
  DFFRX1TF \gr_reg[4][13]  ( .D(N859), .CK(CLK), .RN(RST_N), .Q(N1372) );
  DFFRX1TF \gr_reg[3][13]  ( .D(N867), .CK(CLK), .RN(RST_N), .Q(N1369) );
  DFFRX1TF \gr_reg[2][13]  ( .D(N875), .CK(CLK), .RN(RST_N), .Q(N1366) );
  DFFRX1TF \gr_reg[1][13]  ( .D(N883), .CK(CLK), .RN(RST_N), .Q(N1358) );
  DFFRX1TF \gr_reg[0][13]  ( .D(N891), .CK(CLK), .RN(RST_N), .Q(\GR[0][13] )
         );
  DFFRX1TF \gr_reg[7][15]  ( .D(N833), .CK(CLK), .RN(RST_N), .Q(\GR[7][15] )
         );
  DFFRX1TF \gr_reg[7][14]  ( .D(N834), .CK(CLK), .RN(RST_N), .Q(\GR[7][14] )
         );
  DFFRX1TF \gr_reg[7][12]  ( .D(N836), .CK(CLK), .RN(RST_N), .Q(\GR[7][12] )
         );
  DFFRX1TF \gr_reg[7][11]  ( .D(N837), .CK(CLK), .RN(RST_N), .Q(\GR[7][11] )
         );
  DFFRX1TF \gr_reg[7][10]  ( .D(N838), .CK(CLK), .RN(RST_N), .Q(\GR[7][10] )
         );
  DFFRX1TF \gr_reg[7][9]  ( .D(N839), .CK(CLK), .RN(RST_N), .Q(\GR[7][9] ) );
  DFFRX1TF \gr_reg[7][8]  ( .D(N840), .CK(CLK), .RN(RST_N), .Q(\GR[7][8] ) );
  DFFRX1TF \gr_reg[7][7]  ( .D(N897), .CK(CLK), .RN(RST_N), .Q(\GR[7][7] ) );
  DFFRX1TF \gr_reg[7][6]  ( .D(N898), .CK(CLK), .RN(RST_N), .Q(\GR[7][6] ) );
  DFFRX1TF \gr_reg[7][4]  ( .D(N900), .CK(CLK), .RN(RST_N), .Q(\GR[7][4] ) );
  DFFRX1TF \gr_reg[7][3]  ( .D(N901), .CK(CLK), .RN(RST_N), .Q(\GR[7][3] ) );
  DFFRX1TF \gr_reg[7][2]  ( .D(N902), .CK(CLK), .RN(RST_N), .Q(\GR[7][2] ) );
  DFFRX1TF \gr_reg[7][1]  ( .D(N903), .CK(CLK), .RN(RST_N), .Q(\GR[7][1] ) );
  DFFRX1TF \gr_reg[7][0]  ( .D(N904), .CK(CLK), .RN(RST_N), .Q(\GR[7][0] ) );
  DFFRX1TF \gr_reg[6][15]  ( .D(N841), .CK(CLK), .RN(RST_N), .Q(\GR[6][15] )
         );
  DFFRX1TF \gr_reg[6][14]  ( .D(N842), .CK(CLK), .RN(RST_N), .Q(\GR[6][14] )
         );
  DFFRX1TF \gr_reg[6][12]  ( .D(N844), .CK(CLK), .RN(RST_N), .Q(\GR[6][12] )
         );
  DFFRX1TF \gr_reg[6][11]  ( .D(N845), .CK(CLK), .RN(RST_N), .Q(\GR[6][11] )
         );
  DFFRX1TF \gr_reg[6][10]  ( .D(N846), .CK(CLK), .RN(RST_N), .Q(\GR[6][10] )
         );
  DFFRX1TF \gr_reg[6][9]  ( .D(N847), .CK(CLK), .RN(RST_N), .Q(\GR[6][9] ) );
  DFFRX1TF \gr_reg[6][8]  ( .D(N848), .CK(CLK), .RN(RST_N), .Q(\GR[6][8] ) );
  DFFRX1TF \gr_reg[6][7]  ( .D(N905), .CK(CLK), .RN(RST_N), .Q(\GR[6][7] ) );
  DFFRX1TF \gr_reg[6][6]  ( .D(N906), .CK(CLK), .RN(RST_N), .Q(\GR[6][6] ) );
  DFFRX1TF \gr_reg[6][4]  ( .D(N908), .CK(CLK), .RN(RST_N), .Q(\GR[6][4] ) );
  DFFRX1TF \gr_reg[6][3]  ( .D(N909), .CK(CLK), .RN(RST_N), .Q(\GR[6][3] ) );
  DFFRX1TF \gr_reg[6][2]  ( .D(N910), .CK(CLK), .RN(RST_N), .Q(\GR[6][2] ) );
  DFFRX1TF \gr_reg[6][1]  ( .D(N911), .CK(CLK), .RN(RST_N), .Q(\GR[6][1] ) );
  DFFRX1TF \gr_reg[6][0]  ( .D(N912), .CK(CLK), .RN(RST_N), .Q(\GR[6][0] ) );
  DFFRX1TF \gr_reg[5][15]  ( .D(N849), .CK(CLK), .RN(RST_N), .Q(\GR[5][15] )
         );
  DFFRX1TF \gr_reg[5][14]  ( .D(N850), .CK(CLK), .RN(RST_N), .Q(\GR[5][14] )
         );
  DFFRX1TF \gr_reg[5][12]  ( .D(N852), .CK(CLK), .RN(RST_N), .Q(\GR[5][12] )
         );
  DFFRX1TF \gr_reg[5][11]  ( .D(N853), .CK(CLK), .RN(RST_N), .Q(\GR[5][11] )
         );
  DFFRX1TF \gr_reg[5][10]  ( .D(N854), .CK(CLK), .RN(RST_N), .Q(\GR[5][10] )
         );
  DFFRX1TF \gr_reg[5][9]  ( .D(N855), .CK(CLK), .RN(RST_N), .Q(\GR[5][9] ) );
  DFFRX1TF \gr_reg[5][8]  ( .D(N856), .CK(CLK), .RN(RST_N), .Q(\GR[5][8] ) );
  DFFRX1TF \gr_reg[5][7]  ( .D(N913), .CK(CLK), .RN(RST_N), .Q(\GR[5][7] ) );
  DFFRX1TF \gr_reg[5][6]  ( .D(N914), .CK(CLK), .RN(RST_N), .Q(\GR[5][6] ) );
  DFFRX1TF \gr_reg[5][4]  ( .D(N916), .CK(CLK), .RN(RST_N), .Q(\GR[5][4] ) );
  DFFRX1TF \gr_reg[5][3]  ( .D(N917), .CK(CLK), .RN(RST_N), .Q(\GR[5][3] ) );
  DFFRX1TF \gr_reg[5][2]  ( .D(N918), .CK(CLK), .RN(RST_N), .Q(\GR[5][2] ) );
  DFFRX1TF \gr_reg[5][1]  ( .D(N919), .CK(CLK), .RN(RST_N), .Q(\GR[5][1] ) );
  DFFRX1TF \gr_reg[5][0]  ( .D(N920), .CK(CLK), .RN(RST_N), .Q(\GR[5][0] ) );
  DFFRX1TF \gr_reg[4][15]  ( .D(N857), .CK(CLK), .RN(RST_N), .Q(N1370) );
  DFFRX1TF \gr_reg[4][14]  ( .D(N858), .CK(CLK), .RN(RST_N), .Q(N1371) );
  DFFRX1TF \gr_reg[4][12]  ( .D(N860), .CK(CLK), .RN(RST_N), .Q(N1373) );
  DFFRX1TF \gr_reg[4][11]  ( .D(N861), .CK(CLK), .RN(RST_N), .Q(N1374) );
  DFFRX1TF \gr_reg[4][10]  ( .D(N862), .CK(CLK), .RN(RST_N), .Q(N1375) );
  DFFRX1TF \gr_reg[4][9]  ( .D(N863), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[9])
         );
  DFFRX1TF \gr_reg[4][8]  ( .D(N864), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[8])
         );
  DFFRX1TF \gr_reg[4][7]  ( .D(N921), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[7])
         );
  DFFRX1TF \gr_reg[4][6]  ( .D(N922), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[6])
         );
  DFFRX1TF \gr_reg[4][4]  ( .D(N924), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[4])
         );
  DFFRX1TF \gr_reg[4][3]  ( .D(N925), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[3])
         );
  DFFRX1TF \gr_reg[4][2]  ( .D(N926), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[2])
         );
  DFFRX1TF \gr_reg[4][1]  ( .D(N927), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[1])
         );
  DFFRX1TF \gr_reg[4][0]  ( .D(N928), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[0])
         );
  DFFRX1TF \gr_reg[3][15]  ( .D(N865), .CK(CLK), .RN(RST_N), .Q(N1367) );
  DFFRX1TF \gr_reg[3][14]  ( .D(N866), .CK(CLK), .RN(RST_N), .Q(N1368) );
  DFFRX1TF \gr_reg[3][11]  ( .D(N869), .CK(CLK), .RN(RST_N), .Q(N44), .QN(
        N2070) );
  DFFRX1TF \gr_reg[3][7]  ( .D(N929), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[7])
         );
  DFFRX1TF \gr_reg[3][6]  ( .D(N930), .CK(CLK), .RN(RST_N), .Q(N32), .QN(N193)
         );
  DFFRX1TF \gr_reg[3][4]  ( .D(N932), .CK(CLK), .RN(RST_N), .Q(N39), .QN(N195)
         );
  DFFRX1TF \gr_reg[3][3]  ( .D(N933), .CK(CLK), .RN(RST_N), .Q(N38), .QN(N2010) );
  DFFRX1TF \gr_reg[2][15]  ( .D(N873), .CK(CLK), .RN(RST_N), .Q(N1364) );
  DFFRX1TF \gr_reg[2][14]  ( .D(N874), .CK(CLK), .RN(RST_N), .Q(N1365) );
  DFFRX1TF \gr_reg[2][12]  ( .D(N876), .CK(CLK), .RN(RST_N), .Q(N43), .QN(
        N2050) );
  DFFRX1TF \gr_reg[2][11]  ( .D(N877), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTA[11]) );
  DFFRX1TF \gr_reg[2][10]  ( .D(N878), .CK(CLK), .RN(RST_N), .Q(N42), .QN(N191) );
  DFFRX1TF \gr_reg[2][9]  ( .D(N879), .CK(CLK), .RN(RST_N), .Q(N41), .QN(N290)
         );
  DFFRX1TF \gr_reg[2][8]  ( .D(N880), .CK(CLK), .RN(RST_N), .Q(N40), .QN(N189)
         );
  DFFRX1TF \gr_reg[2][7]  ( .D(N937), .CK(CLK), .RN(RST_N), .Q(N37), .QN(N288)
         );
  DFFRX1TF \gr_reg[2][6]  ( .D(N938), .CK(CLK), .RN(RST_N), .Q(N36), .QN(N2140) );
  DFFRX1TF \gr_reg[2][4]  ( .D(N940), .CK(CLK), .RN(RST_N), .Q(N35), .QN(N286)
         );
  DFFRX1TF \gr_reg[2][3]  ( .D(N941), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[3])
         );
  DFFRX1TF \gr_reg[2][2]  ( .D(N942), .CK(CLK), .RN(RST_N), .Q(N34), .QN(N218)
         );
  DFFRX1TF \gr_reg[2][1]  ( .D(N943), .CK(CLK), .RN(RST_N), .Q(N33), .QN(N2030) );
  DFFRX1TF \gr_reg[1][15]  ( .D(N881), .CK(CLK), .RN(RST_N), .Q(N1356) );
  DFFRX1TF \gr_reg[1][14]  ( .D(N882), .CK(CLK), .RN(RST_N), .Q(N1357) );
  DFFRX1TF \gr_reg[1][12]  ( .D(N884), .CK(CLK), .RN(RST_N), .Q(N1359) );
  DFFRX1TF \gr_reg[1][11]  ( .D(N885), .CK(CLK), .RN(RST_N), .Q(N1360) );
  DFFRX1TF \gr_reg[1][10]  ( .D(N886), .CK(CLK), .RN(RST_N), .Q(N1361) );
  DFFRX1TF \gr_reg[1][9]  ( .D(N887), .CK(CLK), .RN(RST_N), .Q(N1362) );
  DFFRX1TF \gr_reg[1][8]  ( .D(N888), .CK(CLK), .RN(RST_N), .Q(N1363) );
  DFFRX1TF \gr_reg[1][6]  ( .D(N946), .CK(CLK), .RN(RST_N), .Q(\IO_CONTROL[6] ) );
  DFFRX1TF \gr_reg[1][1]  ( .D(N951), .CK(CLK), .RN(RST_N), .Q(\IO_CONTROL[1] ) );
  DFFRX1TF \gr_reg[1][0]  ( .D(N952), .CK(CLK), .RN(RST_N), .Q(\IO_CONTROL[0] ) );
  DFFRX1TF \gr_reg[0][15]  ( .D(N889), .CK(CLK), .RN(RST_N), .Q(\GR[0][15] )
         );
  DFFRX1TF \gr_reg[0][14]  ( .D(N890), .CK(CLK), .RN(RST_N), .Q(\GR[0][14] )
         );
  DFFRX1TF \gr_reg[0][12]  ( .D(N892), .CK(CLK), .RN(RST_N), .Q(\GR[0][12] )
         );
  DFFRX1TF \gr_reg[0][11]  ( .D(N893), .CK(CLK), .RN(RST_N), .Q(\GR[0][11] )
         );
  DFFRX1TF \gr_reg[0][10]  ( .D(N894), .CK(CLK), .RN(RST_N), .Q(\GR[0][10] )
         );
  DFFRX1TF \gr_reg[0][9]  ( .D(N895), .CK(CLK), .RN(RST_N), .Q(\GR[0][9] ) );
  DFFRX1TF \gr_reg[0][8]  ( .D(N896), .CK(CLK), .RN(RST_N), .Q(\GR[0][8] ) );
  DFFRX1TF \gr_reg[0][7]  ( .D(N953), .CK(CLK), .RN(RST_N), .Q(\GR[0][7] ) );
  DFFRX1TF \gr_reg[0][6]  ( .D(N954), .CK(CLK), .RN(RST_N), .Q(\GR[0][6] ) );
  DFFRX1TF \gr_reg[0][4]  ( .D(N956), .CK(CLK), .RN(RST_N), .Q(\GR[0][4] ) );
  DFFRX1TF \gr_reg[0][3]  ( .D(N957), .CK(CLK), .RN(RST_N), .Q(\GR[0][3] ) );
  DFFRX1TF \gr_reg[0][2]  ( .D(N958), .CK(CLK), .RN(RST_N), .Q(\GR[0][2] ) );
  DFFRX1TF \gr_reg[0][1]  ( .D(N959), .CK(CLK), .RN(RST_N), .Q(\GR[0][1] ) );
  DFFRX1TF \gr_reg[0][0]  ( .D(N960), .CK(CLK), .RN(RST_N), .Q(\GR[0][0] ) );
  DFFRX1TF \gr_reg[7][5]  ( .D(N899), .CK(CLK), .RN(RST_N), .Q(\GR[7][5] ) );
  DFFRX1TF \gr_reg[6][5]  ( .D(N907), .CK(CLK), .RN(RST_N), .Q(\GR[6][5] ) );
  DFFRX1TF \gr_reg[5][5]  ( .D(N915), .CK(CLK), .RN(RST_N), .Q(\GR[5][5] ) );
  DFFRX1TF \gr_reg[4][5]  ( .D(N923), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[5])
         );
  DFFRX1TF \gr_reg[3][5]  ( .D(N931), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[5])
         );
  DFFRX1TF \gr_reg[2][5]  ( .D(N939), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[5])
         );
  DFFRX1TF \gr_reg[1][5]  ( .D(N947), .CK(CLK), .RN(RST_N), .Q(\IO_CONTROL[5] ), .QN(\IO_CONTROL[5]_BAR ) );
  DFFRX1TF \gr_reg[0][5]  ( .D(N955), .CK(CLK), .RN(RST_N), .Q(\GR[0][5] ) );
  DFFNSRX2TF lowest_bit_reg ( .D(N962), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        I_ADDR[0]), .QN(N347) );
  DFFRX2TF \gr_reg[3][9]  ( .D(N871), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[9])
         );
  DFFRX2TF \gr_reg[3][1]  ( .D(N935), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[1])
         );
  DFFRX2TF \gr_reg[3][12]  ( .D(N868), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTB[12]) );
  DFFRX2TF \gr_reg[2][0]  ( .D(N944), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[0])
         );
  DFFRX2TF \gr_reg[3][0]  ( .D(N936), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[0])
         );
  DFFRX2TF \gr_reg[3][2]  ( .D(N934), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[2])
         );
  DFFRX2TF \gr_reg[1][4]  ( .D(N948), .CK(CLK), .RN(RST_N), .Q(\IO_CONTROL[4] ) );
  DFFRX2TF \gr_reg[3][10]  ( .D(N870), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTB[10]) );
  DFFRX2TF \gr_reg[1][7]  ( .D(N945), .CK(CLK), .RN(RST_N), .Q(\IO_CONTROL[7] ) );
  DFFRX2TF \gr_reg[1][2]  ( .D(N950), .CK(CLK), .RN(RST_N), .Q(\IO_CONTROL[2] ) );
  DFFNSRX2TF \reg_C_reg[8]  ( .D(N440), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[9]) );
  DFFRX2TF \gr_reg[3][8]  ( .D(N872), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[8])
         );
  DFFRX2TF \gr_reg[1][3]  ( .D(N949), .CK(CLK), .RN(RST_N), .Q(\IO_CONTROL[3] ) );
  DFFRX2TF \reg_B_reg[1]  ( .D(N473), .CK(CLK), .RN(RST_N), .Q(REG_B[1]), .QN(
        N355) );
  DFFRX2TF \id_ir_reg[15]  ( .D(N517), .CK(CLK), .RN(RST_N), .Q(N29), .QN(N358) );
  DFFRX2TF \reg_B_reg[0]  ( .D(N474), .CK(CLK), .RN(RST_N), .Q(REG_B[0]), .QN(
        N354) );
  DFFRX2TF \id_ir_reg[13]  ( .D(N519), .CK(CLK), .RN(RST_N), .Q(CODE_TYPE[2]), 
        .QN(N346) );
  NOR4X4TF U3 ( .A(STATE[3]), .B(N552), .C(STATE[1]), .D(N348), .Y(N1104) );
  NOR3X1TF U4 ( .A(CODE_TYPE[3]), .B(N2110), .C(N1103), .Y(N1088) );
  INVX2TF U5 ( .A(N376), .Y(N1044) );
  NAND3X1TF U6 ( .A(N2000), .B(N634), .C(N306), .Y(N1064) );
  AOI2BB2X1TF U7 ( .B0(N1010), .B1(N604), .A0N(N1015), .A1N(N979), .Y(N1) );
  AOI22X1TF U8 ( .A0(REG_A[7]), .A1(N608), .B0(N387), .B1(N343), .Y(N2) );
  AOI32X1TF U9 ( .A0(N376), .A1(N1), .A2(N2), .B0(N580), .B1(N1), .Y(N3) );
  AO21X1TF U10 ( .A0(N580), .A1(N386), .B0(N1047), .Y(N4) );
  AOI22X1TF U11 ( .A0(REG_A[7]), .A1(N4), .B0(N612), .B1(N1011), .Y(N5) );
  AOI22X1TF U12 ( .A0(N988), .A1(N978), .B0(N490), .B1(N268), .Y(N6) );
  OAI211X1TF U13 ( .A0(N992), .A1(N1017), .B0(N5), .C0(N6), .Y(N7) );
  AOI211X1TF U14 ( .A0(N546), .A1(N456), .B0(N3), .C0(N7), .Y(N592) );
  NOR2BX1TF U15 ( .AN(N1102), .B(N359), .Y(N1099) );
  NAND3BX1TF U16 ( .AN(CODE_TYPE[3]), .B(N648), .C(N2000), .Y(N647) );
  AOI21X1TF U17 ( .A0(REG_A[5]), .A1(N2130), .B0(N764), .Y(N8) );
  NAND3X1TF U18 ( .A(N812), .B(N774), .C(N8), .Y(N1011) );
  AO22X1TF U19 ( .A0(REG_A[8]), .A1(N292), .B0(N386), .B1(N341), .Y(N9) );
  NOR2X1TF U20 ( .A(N1044), .B(N9), .Y(N10) );
  AOI22X1TF U21 ( .A0(N612), .A1(N985), .B0(N984), .B1(N604), .Y(N11) );
  OAI21X1TF U22 ( .A0(N986), .A1(N992), .B0(N11), .Y(N12) );
  AOI21X1TF U23 ( .A0(N579), .A1(N388), .B0(N1047), .Y(N13) );
  OAI22X1TF U24 ( .A0(N341), .A1(N13), .B0(N983), .B1(N982), .Y(N14) );
  AOI211X1TF U25 ( .A0(N378), .A1(N457), .B0(N12), .C0(N14), .Y(N15) );
  AOI22X1TF U26 ( .A0(N988), .A1(N987), .B0(N491), .B1(N267), .Y(N16) );
  OAI211X1TF U27 ( .A0(N579), .A1(N10), .B0(N15), .C0(N16), .Y(N1055) );
  OA21XLTF U28 ( .A0(I_ADDR[1]), .A1(I_ADDR[2]), .B0(N699), .Y(N17) );
  AOI222XLTF U29 ( .A0(I_ADDR[2]), .A1(N711), .B0(N719), .B1(D_ADDR[2]), .C0(
        N709), .C1(N17), .Y(N726) );
  OAI211X1TF U30 ( .A0(N30), .A1(N362), .B0(N789), .C0(N759), .Y(N18) );
  NOR2X1TF U31 ( .A(N758), .B(N18), .Y(N1037) );
  AOI211X1TF U32 ( .A0(REG_A[11]), .A1(N302), .B0(N769), .C0(N763), .Y(N19) );
  NAND2X1TF U33 ( .A(N811), .B(N19), .Y(N1012) );
  AOI2BB1X1TF U34 ( .A0N(N1068), .A1N(N1069), .B0(N1052), .Y(N589) );
  OA21XLTF U35 ( .A0(N710), .A1(I_ADDR[7]), .B0(N715), .Y(N20) );
  AOI222XLTF U36 ( .A0(I_ADDR[7]), .A1(N711), .B0(N719), .B1(D_ADDR[7]), .C0(
        N709), .C1(N20), .Y(N721) );
  NOR3X1TF U37 ( .A(N601), .B(N268), .C(N292), .Y(N21) );
  NAND3X1TF U38 ( .A(N632), .B(N357), .C(N21), .Y(N567) );
  NAND3BX1TF U39 ( .AN(N91), .B(N89), .C(N90), .Y(N1147) );
  NAND3BX1TF U40 ( .AN(N94), .B(N92), .C(N93), .Y(N1219) );
  NAND3BX1TF U41 ( .AN(N97), .B(N95), .C(N96), .Y(N1291) );
  AOI21X1TF U42 ( .A0(N1064), .A1(N359), .B0(N29), .Y(N22) );
  NAND3X1TF U43 ( .A(N1104), .B(N1086), .C(N22), .Y(N220) );
  NOR4BBX1TF U44 ( .AN(N593), .BN(N589), .C(N1059), .D(N1058), .Y(N23) );
  NAND4BX1TF U45 ( .AN(N1061), .B(N23), .C(N594), .D(N592), .Y(N24) );
  NOR4XLTF U46 ( .A(N1056), .B(N1057), .C(N1060), .D(N24), .Y(N25) );
  NAND4BX1TF U47 ( .AN(N1055), .B(N588), .C(N25), .D(N600), .Y(N26) );
  NAND4X1TF U48 ( .A(N576), .B(N590), .C(N598), .D(N585), .Y(N27) );
  OAI22X1TF U49 ( .A0(N589), .A1(N368), .B0(N26), .B1(N27), .Y(N4570) );
  AOI21X1TF U50 ( .A0(N699), .A1(N373), .B0(N713), .Y(N28) );
  AOI222XLTF U51 ( .A0(I_ADDR[3]), .A1(N711), .B0(N28), .B1(N700), .C0(N719), 
        .C1(D_ADDR[3]), .Y(N725) );
  INVX2TF U52 ( .A(CODE_TYPE[2]), .Y(N1990) );
  INVX2TF U53 ( .A(REG_B[0]), .Y(N197) );
  NAND2X2TF U54 ( .A(REG_B[1]), .B(N354), .Y(N30) );
  AO22X1TF U55 ( .A0(N1138), .A1(N1137), .B0(N5670), .B1(N1139), .Y(N31) );
  AOI22XLTF U56 ( .A0(N379), .A1(\IO_CONTROL[2] ), .B0(N2540), .B1(
        IO_DATAOUTB[2]), .Y(N1157) );
  AOI22XLTF U57 ( .A0(N277), .A1(\IO_CONTROL[2] ), .B0(N2520), .B1(
        IO_DATAOUTB[2]), .Y(N1229) );
  AOI22XLTF U58 ( .A0(N280), .A1(\IO_CONTROL[2] ), .B0(N256), .B1(
        IO_DATAOUTB[2]), .Y(N1301) );
  NAND2BX4TF U59 ( .AN(REG_A[0]), .B(REG_B[0]), .Y(SUB_X_300_4_N16) );
  CLKINVX1TF U67 ( .A(N1086), .Y(N1087) );
  OAI2BB1X1TF U68 ( .A0N(N396), .A1N(N611), .B0(N395), .Y(N1028) );
  NOR2X1TF U69 ( .A(N1064), .B(N390), .Y(N609) );
  OR3X1TF U70 ( .A(N97), .B(N95), .C(N352), .Y(N1285) );
  OR3X1TF U71 ( .A(N94), .B(N92), .C(N93), .Y(N1212) );
  OR3X1TF U72 ( .A(N91), .B(N89), .C(N351), .Y(N1141) );
  OAI211X2TF U73 ( .A0(N557), .A1(N350), .B0(N556), .C0(N555), .Y(N558) );
  OAI2BB2XLTF U74 ( .B0(N575), .B1(N630), .A0N(N404), .A1N(N612), .Y(N405) );
  OAI2BB2XLTF U75 ( .B0(N439), .B1(N582), .A0N(N454), .A1N(N378), .Y(N441) );
  INVX1TF U76 ( .A(N827), .Y(N828) );
  OR2X2TF U77 ( .A(N661), .B(N681), .Y(N656) );
  CLKINVX2TF U78 ( .A(N996), .Y(N528) );
  OR2X2TF U79 ( .A(N659), .B(N684), .Y(N657) );
  OR2X2TF U80 ( .A(N689), .B(N688), .Y(N698) );
  OR2X2TF U81 ( .A(N661), .B(N684), .Y(N658) );
  OR2X2TF U82 ( .A(N684), .B(N686), .Y(N683) );
  OR2X2TF U83 ( .A(N659), .B(N689), .Y(N660) );
  OR2X2TF U84 ( .A(N681), .B(N688), .Y(N682) );
  OR2X2TF U85 ( .A(N678), .B(N659), .Y(N652) );
  OR2X2TF U86 ( .A(N681), .B(N686), .Y(N680) );
  OR2X2TF U87 ( .A(N678), .B(N688), .Y(N679) );
  OR2X2TF U88 ( .A(N661), .B(N689), .Y(N670) );
  OR2X2TF U89 ( .A(N678), .B(N686), .Y(N676) );
  AOI22X1TF U90 ( .A0(N305), .A1(N167), .B0(N304), .B1(N204), .Y(N1115) );
  AOI22X1TF U91 ( .A0(N305), .A1(N164), .B0(N304), .B1(N201), .Y(N1112) );
  AOI22X1TF U92 ( .A0(N305), .A1(N162), .B0(N304), .B1(N199), .Y(N1110) );
  AOI22X1TF U93 ( .A0(N305), .A1(N172), .B0(N304), .B1(N209), .Y(N1120) );
  AOI22X1TF U94 ( .A0(N1126), .A1(N177), .B0(N1125), .B1(N214), .Y(N1127) );
  AOI22X1TF U95 ( .A0(N1126), .A1(N173), .B0(N1125), .B1(N210), .Y(N1121) );
  AOI22X1TF U96 ( .A0(N1126), .A1(N171), .B0(N1125), .B1(N208), .Y(N1119) );
  AOI22X1TF U97 ( .A0(N1126), .A1(N176), .B0(N1125), .B1(N213), .Y(N1124) );
  AOI22X1TF U98 ( .A0(N305), .A1(N165), .B0(N304), .B1(N202), .Y(N1113) );
  AOI22X1TF U99 ( .A0(N1126), .A1(N163), .B0(N1125), .B1(N200), .Y(N1111) );
  AOI22X1TF U100 ( .A0(N1126), .A1(N166), .B0(N1125), .B1(N203), .Y(N1114) );
  AOI22X1TF U101 ( .A0(N1126), .A1(N169), .B0(N1125), .B1(N206), .Y(N1117) );
  AOI22X1TF U102 ( .A0(N1126), .A1(N175), .B0(N1125), .B1(N212), .Y(N1123) );
  AOI22X1TF U103 ( .A0(N1126), .A1(N170), .B0(N1125), .B1(N207), .Y(N1118) );
  AOI22X1TF U104 ( .A0(N305), .A1(N168), .B0(N304), .B1(N205), .Y(N1116) );
  AOI22X1TF U105 ( .A0(N1126), .A1(N174), .B0(N1125), .B1(N211), .Y(N1122) );
  INVX2TF U106 ( .A(N1132), .Y(N264) );
  OAI211X1TF U107 ( .A0(N1130), .A1(N1107), .B0(N1108), .C0(N1109), .Y(N1128)
         );
  NAND4BXLTF U108 ( .AN(N158), .B(N737), .C(N736), .D(N735), .Y(NEXT_STATE[3])
         );
  OR2X2TF U109 ( .A(N1130), .B(N1129), .Y(N1132) );
  OAI211X1TF U110 ( .A0(STATE[3]), .A1(N645), .B0(N644), .C0(N735), .Y(N962)
         );
  CLKINVX2TF U111 ( .A(N671), .Y(N303) );
  AOI22X1TF U112 ( .A0(N282), .A1(\GR[0][2] ), .B0(N258), .B1(N34), .Y(N1156)
         );
  NAND2XLTF U113 ( .A(N1031), .B(REG_A[10]), .Y(N753) );
  AOI22X1TF U114 ( .A0(N284), .A1(\GR[0][2] ), .B0(N262), .B1(N34), .Y(N1300)
         );
  AOI22X1TF U115 ( .A0(N1143), .A1(IO_OFFSET[3]), .B0(N269), .B1(\GR[6][3] ), 
        .Y(N1162) );
  AOI22X1TF U116 ( .A0(N1287), .A1(IO_OFFSET[0]), .B0(N271), .B1(\GR[6][0] ), 
        .Y(N1294) );
  AOI22X1TF U117 ( .A0(N1143), .A1(N1371), .B0(N269), .B1(\GR[6][14] ), .Y(
        N1206) );
  AOI22X1TF U118 ( .A0(N1143), .A1(N1374), .B0(N269), .B1(\GR[6][11] ), .Y(
        N1194) );
  AOI22X1TF U119 ( .A0(N1215), .A1(N1371), .B0(N273), .B1(\GR[6][14] ), .Y(
        N1278) );
  AOI22X1TF U120 ( .A0(N1287), .A1(N1373), .B0(N271), .B1(\GR[6][12] ), .Y(
        N1342) );
  AOI22X1TF U121 ( .A0(N226), .A1(\GR[0][2] ), .B0(N275), .B1(N34), .Y(N1228)
         );
  NAND4XLTF U122 ( .A(N734), .B(N732), .C(N731), .D(N730), .Y(NEXT_STATE[1])
         );
  AOI22X1TF U123 ( .A0(N226), .A1(\GR[0][8] ), .B0(N275), .B1(N40), .Y(N1252)
         );
  AOI22X1TF U124 ( .A0(N1287), .A1(IO_OFFSET[9]), .B0(N271), .B1(\GR[6][9] ), 
        .Y(N1330) );
  AOI22X1TF U125 ( .A0(N1287), .A1(IO_OFFSET[2]), .B0(N271), .B1(\GR[6][2] ), 
        .Y(N1302) );
  AOI22X1TF U126 ( .A0(N226), .A1(\GR[0][1] ), .B0(N275), .B1(N33), .Y(N1224)
         );
  AOI22X1TF U127 ( .A0(N1215), .A1(IO_OFFSET[1]), .B0(N273), .B1(\GR[6][1] ), 
        .Y(N1226) );
  AOI22X1TF U128 ( .A0(N226), .A1(\GR[0][6] ), .B0(N275), .B1(N36), .Y(N1244)
         );
  AOI22X1TF U129 ( .A0(N1215), .A1(IO_OFFSET[3]), .B0(N273), .B1(\GR[6][3] ), 
        .Y(N1234) );
  AOI22X1TF U130 ( .A0(N1287), .A1(IO_OFFSET[1]), .B0(N271), .B1(\GR[6][1] ), 
        .Y(N1298) );
  AOI22X1TF U131 ( .A0(N1215), .A1(IO_OFFSET[0]), .B0(N273), .B1(\GR[6][0] ), 
        .Y(N1222) );
  AOI22X1TF U132 ( .A0(N1287), .A1(IO_OFFSET[3]), .B0(N271), .B1(\GR[6][3] ), 
        .Y(N1306) );
  AOI22X1TF U133 ( .A0(N1143), .A1(IO_OFFSET[1]), .B0(N269), .B1(\GR[6][1] ), 
        .Y(N1154) );
  AOI22X1TF U134 ( .A0(N1215), .A1(N1374), .B0(N273), .B1(\GR[6][11] ), .Y(
        N1266) );
  AOI22X1TF U135 ( .A0(N1143), .A1(IO_OFFSET[8]), .B0(N269), .B1(\GR[6][8] ), 
        .Y(N1182) );
  AOI22X1TF U136 ( .A0(N1143), .A1(IO_OFFSET[6]), .B0(N269), .B1(\GR[6][6] ), 
        .Y(N1174) );
  AOI22X1TF U137 ( .A0(N1215), .A1(IO_OFFSET[8]), .B0(N273), .B1(\GR[6][8] ), 
        .Y(N1254) );
  NOR2X4TF U138 ( .A(STATE[2]), .B(N732), .Y(N651) );
  NAND2XLTF U139 ( .A(N2000), .B(N306), .Y(N1066) );
  NOR2X4TF U140 ( .A(N198), .B(REG_B[1]), .Y(N1031) );
  NAND4XLTF U141 ( .A(I_ADDR[0]), .B(N643), .C(N737), .D(N1130), .Y(N644) );
  NAND2X2TF U142 ( .A(N198), .B(N355), .Y(N756) );
  AND2X2TF U143 ( .A(N198), .B(REG_B[1]), .Y(N808) );
  NOR2X4TF U144 ( .A(N732), .B(N348), .Y(N650) );
  NAND2XLTF U145 ( .A(N307), .B(N346), .Y(N1065) );
  OR3X1TF U146 ( .A(N91), .B(N89), .C(N90), .Y(N1140) );
  OR3X1TF U147 ( .A(N89), .B(N335), .C(N351), .Y(N1144) );
  OR3X1TF U148 ( .A(N94), .B(N92), .C(N353), .Y(N1213) );
  OR3X1TF U149 ( .A(N94), .B(N93), .C(N371), .Y(N1214) );
  OR3X1TF U150 ( .A(N92), .B(N337), .C(N353), .Y(N1216) );
  OR3X1TF U151 ( .A(N95), .B(N336), .C(N352), .Y(N1288) );
  OR3X1TF U152 ( .A(N97), .B(N96), .C(N370), .Y(N1286) );
  OR3X1TF U153 ( .A(N97), .B(N95), .C(N96), .Y(N1284) );
  INVX2TF U154 ( .A(N189), .Y(IO_DATAOUTA[8]) );
  INVX2TF U155 ( .A(N191), .Y(IO_DATAOUTA[10]) );
  INVX2TF U156 ( .A(N193), .Y(IO_DATAOUTB[6]) );
  INVX2TF U157 ( .A(N195), .Y(IO_DATAOUTB[4]) );
  INVX2TF U158 ( .A(N197), .Y(N198) );
  INVX2TF U159 ( .A(N1990), .Y(N2000) );
  INVX2TF U160 ( .A(N2010), .Y(IO_DATAOUTB[3]) );
  INVX2TF U161 ( .A(N2030), .Y(IO_DATAOUTA[1]) );
  INVX2TF U162 ( .A(N2050), .Y(IO_DATAOUTA[12]) );
  INVX2TF U163 ( .A(N2070), .Y(IO_DATAOUTB[11]) );
  INVX2TF U164 ( .A(N808), .Y(N2090) );
  INVX2TF U165 ( .A(N808), .Y(N2100) );
  INVX2TF U166 ( .A(N358), .Y(N2110) );
  INVX2TF U167 ( .A(N1030), .Y(N2120) );
  INVX2TF U168 ( .A(N2120), .Y(N2130) );
  INVX2TF U169 ( .A(N2140), .Y(IO_DATAOUTA[6]) );
  INVX2TF U170 ( .A(N597), .Y(N216) );
  INVX2TF U171 ( .A(N216), .Y(N217) );
  INVX2TF U172 ( .A(N218), .Y(IO_DATAOUTA[2]) );
  INVX2TF U173 ( .A(N220), .Y(N221) );
  INVX2TF U174 ( .A(N220), .Y(N222) );
  INVX2TF U175 ( .A(N1128), .Y(N223) );
  INVX2TF U176 ( .A(N223), .Y(N224) );
  INVX2TF U177 ( .A(N223), .Y(N225) );
  INVX2TF U178 ( .A(N1212), .Y(N226) );
  INVX2TF U179 ( .A(N1212), .Y(N227) );
  INVX2TF U180 ( .A(N680), .Y(N228) );
  INVX2TF U181 ( .A(N680), .Y(N229) );
  INVX2TF U182 ( .A(N698), .Y(N230) );
  INVX2TF U183 ( .A(N698), .Y(N231) );
  INVX2TF U184 ( .A(N679), .Y(N232) );
  INVX2TF U185 ( .A(N679), .Y(N233) );
  INVX2TF U186 ( .A(N682), .Y(N234) );
  INVX2TF U187 ( .A(N682), .Y(N235) );
  INVX2TF U188 ( .A(N683), .Y(N236) );
  INVX2TF U189 ( .A(N683), .Y(N237) );
  INVX2TF U190 ( .A(N676), .Y(N238) );
  INVX2TF U191 ( .A(N676), .Y(N2390) );
  INVX2TF U192 ( .A(N657), .Y(N2400) );
  INVX2TF U193 ( .A(N657), .Y(N2410) );
  INVX2TF U194 ( .A(N656), .Y(N2420) );
  INVX2TF U195 ( .A(N656), .Y(N2430) );
  INVX2TF U196 ( .A(N670), .Y(N2440) );
  INVX2TF U197 ( .A(N670), .Y(N2450) );
  INVX2TF U198 ( .A(N652), .Y(N2460) );
  INVX2TF U199 ( .A(N652), .Y(N2470) );
  INVX2TF U200 ( .A(N658), .Y(N2480) );
  INVX2TF U201 ( .A(N658), .Y(N2490) );
  INVX2TF U202 ( .A(N660), .Y(N2500) );
  INVX2TF U203 ( .A(N660), .Y(N2510) );
  INVX2TF U204 ( .A(N1219), .Y(N2520) );
  INVX2TF U205 ( .A(N1219), .Y(N2530) );
  INVX2TF U206 ( .A(N1147), .Y(N2540) );
  INVX2TF U207 ( .A(N1147), .Y(N255) );
  INVX2TF U208 ( .A(N1291), .Y(N256) );
  INVX2TF U209 ( .A(N1291), .Y(N257) );
  INVX2TF U210 ( .A(N1141), .Y(N258) );
  INVX2TF U211 ( .A(N1141), .Y(N261) );
  INVX2TF U212 ( .A(N1285), .Y(N262) );
  INVX2TF U213 ( .A(N1285), .Y(N263) );
  INVX2TF U214 ( .A(N1132), .Y(N265) );
  INVX2TF U215 ( .A(N1028), .Y(N266) );
  INVX2TF U216 ( .A(N266), .Y(N267) );
  INVX2TF U217 ( .A(N266), .Y(N268) );
  OAI31X4TF U218 ( .A0(N1088), .A1(N1106), .A2(N1087), .B0(N1104), .Y(N1094)
         );
  NOR2X2TF U219 ( .A(N640), .B(N671), .Y(N709) );
  AOI211X1TF U220 ( .A0(N1063), .A1(N610), .B0(N1047), .C0(N609), .Y(N632) );
  NOR2BX2TF U221 ( .AN(N29), .B(CODE_TYPE[3]), .Y(N610) );
  INVX2TF U222 ( .A(N1144), .Y(N269) );
  INVX2TF U223 ( .A(N1144), .Y(N270) );
  INVX2TF U224 ( .A(N1288), .Y(N271) );
  INVX2TF U225 ( .A(N1288), .Y(N272) );
  INVX2TF U226 ( .A(N1216), .Y(N273) );
  INVX2TF U227 ( .A(N1216), .Y(N274) );
  INVX2TF U228 ( .A(N1213), .Y(N275) );
  INVX2TF U229 ( .A(N1213), .Y(N276) );
  INVX2TF U230 ( .A(N1214), .Y(N277) );
  INVX2TF U231 ( .A(N1214), .Y(N278) );
  INVX2TF U232 ( .A(N1286), .Y(N280) );
  INVX2TF U233 ( .A(N1286), .Y(N281) );
  AOI22XLTF U234 ( .A0(N226), .A1(\GR[0][0] ), .B0(N275), .B1(IO_DATAOUTA[0]), 
        .Y(N1220) );
  AOI22XLTF U235 ( .A0(N226), .A1(\GR[0][5] ), .B0(N275), .B1(IO_DATAOUTA[5]), 
        .Y(N1240) );
  INVX2TF U236 ( .A(N1140), .Y(N282) );
  INVX2TF U237 ( .A(N1140), .Y(N283) );
  INVX2TF U238 ( .A(N1284), .Y(N284) );
  INVX2TF U239 ( .A(N1284), .Y(N285) );
  INVX2TF U240 ( .A(N286), .Y(IO_DATAOUTA[4]) );
  INVX2TF U241 ( .A(N288), .Y(IO_DATAOUTA[7]) );
  INVX2TF U242 ( .A(N290), .Y(IO_DATAOUTA[9]) );
  INVX2TF U243 ( .A(N1013), .Y(N292) );
  CLKBUFX2TF U244 ( .A(N596), .Y(N293) );
  NOR2X1TF U245 ( .A(N415), .B(N1064), .Y(N596) );
  CLKBUFX2TF U246 ( .A(N687), .Y(N294) );
  NOR2X2TF U247 ( .A(N689), .B(N686), .Y(N687) );
  CLKBUFX2TF U248 ( .A(N685), .Y(N295) );
  NOR2X2TF U249 ( .A(N684), .B(N688), .Y(N685) );
  CLKBUFX2TF U250 ( .A(N654), .Y(N296) );
  NOR2X2TF U251 ( .A(N678), .B(N661), .Y(N654) );
  CLKBUFX2TF U252 ( .A(N655), .Y(N297) );
  NOR2X2TF U253 ( .A(N659), .B(N681), .Y(N655) );
  CLKBUFX2TF U254 ( .A(N379), .Y(N298) );
  CLKBUFX2TF U255 ( .A(N1142), .Y(N379) );
  CLKBUFX2TF U256 ( .A(N380), .Y(N299) );
  CLKBUFX2TF U257 ( .A(N1145), .Y(N380) );
  CLKBUFX2TF U258 ( .A(N384), .Y(N300) );
  CLKBUFX2TF U259 ( .A(N1289), .Y(N384) );
  CLKBUFX2TF U260 ( .A(N382), .Y(N301) );
  CLKBUFX2TF U261 ( .A(N1217), .Y(N382) );
  INVX2TF U262 ( .A(N762), .Y(N302) );
  AOI22XLTF U263 ( .A0(REG_B[2]), .A1(N971), .B0(N967), .B1(N356), .Y(N751) );
  INVX2TF U264 ( .A(N1109), .Y(N304) );
  INVX2TF U265 ( .A(N1108), .Y(N305) );
  NOR2X2TF U266 ( .A(REG_B[3]), .B(N356), .Y(N1043) );
  NOR2X2TF U267 ( .A(STATE[3]), .B(STATE[2]), .Y(N1135) );
  AOI211X2TF U268 ( .A0(N1063), .A1(N29), .B0(N607), .C0(N1099), .Y(N1086) );
  INVX2TF U269 ( .A(N306), .Y(N307) );
  NAND2X1TF U270 ( .A(N634), .B(CODE_TYPE[1]), .Y(N648) );
  NAND2X1TF U271 ( .A(N615), .B(CODE_TYPE[1]), .Y(N761) );
  NAND2X1TF U272 ( .A(CODE_TYPE[1]), .B(N1088), .Y(N972) );
  CLKBUFX2TF U273 ( .A(N1143), .Y(N308) );
  CLKBUFX2TF U274 ( .A(N1287), .Y(N309) );
  CLKBUFX2TF U275 ( .A(N1215), .Y(N310) );
  XOR2X1TF U276 ( .A(REG_A[0]), .B(N198), .Y(N483) );
  CMPR32X2TF U277 ( .A(N355), .B(REG_A[1]), .C(SUB_X_300_4_N16), .CO(
        SUB_X_300_4_N15), .S(N484) );
  INVX2TF U278 ( .A(SUB_X_300_4_N1), .Y(N499) );
  ADDFHX4TF U279 ( .A(N572), .B(REG_A[15]), .CI(SUB_X_300_4_N2), .CO(
        SUB_X_300_4_N1), .S(N498) );
  NAND2X2TF U280 ( .A(N464), .B(N546), .Y(N556) );
  XOR2X4TF U281 ( .A(N588), .B(N560), .Y(N565) );
  XOR2X2TF U282 ( .A(N600), .B(N559), .Y(N560) );
  XOR2X4TF U283 ( .A(N598), .B(N1060), .Y(N559) );
  OAI21X4TF U284 ( .A0(N565), .A1(N1053), .B0(N564), .Y(N424) );
  AO21X1TF U285 ( .A0(IO_DATAINA[3]), .A1(N597), .B0(N569), .Y(N430) );
  CLKBUFX2TF U286 ( .A(N546), .Y(N378) );
  OAI22XLTF U287 ( .A0(N29), .A1(N1103), .B0(N1102), .B1(N1101), .Y(N1105) );
  AOI21X4TF U288 ( .A0(N498), .A1(N268), .B0(N558), .Y(N588) );
  AO21X1TF U289 ( .A0(IO_DATAINA[4]), .A1(N597), .B0(N584), .Y(N432) );
  INVX2TF U290 ( .A(N968), .Y(N612) );
  NAND2X2TF U291 ( .A(N5670), .B(CODE_TYPE[2]), .Y(N1103) );
  NAND2X1TF U292 ( .A(N603), .B(N610), .Y(N415) );
  CLKBUFX2TF U293 ( .A(N1052), .Y(N377) );
  AOI211X1TF U294 ( .A0(N1010), .A1(N612), .B0(N821), .C0(N543), .Y(N576) );
  OAI211X1TF U295 ( .A0(N1039), .A1(N968), .B0(N801), .C0(N422), .Y(N1058) );
  AOI31XLTF U296 ( .A0(N1102), .A1(N633), .A2(N306), .B0(N736), .Y(N159) );
  NAND2X1TF U297 ( .A(N5670), .B(N1106), .Y(N672) );
  NAND2X2TF U298 ( .A(N611), .B(N1063), .Y(N357) );
  OAI21X1TF U299 ( .A0(STATE[1]), .A1(N631), .B0(N671), .Y(N157) );
  NAND2X1TF U300 ( .A(N677), .B(N369), .Y(N686) );
  NAND2X1TF U301 ( .A(N89), .B(N677), .Y(N688) );
  NAND2X1TF U302 ( .A(N89), .B(N653), .Y(N661) );
  NAND2X1TF U303 ( .A(N369), .B(N653), .Y(N659) );
  AOI32X1TF U304 ( .A0(N611), .A1(N672), .A2(N1103), .B0(N649), .B1(N672), .Y(
        N673) );
  NOR4X1TF U305 ( .A(CODE_TYPE[3]), .B(N29), .C(N2000), .D(N306), .Y(N1106) );
  NAND2X1TF U306 ( .A(STATE[3]), .B(N1136), .Y(N732) );
  NOR2X1TF U307 ( .A(N552), .B(N375), .Y(N1136) );
  CLKBUFX6TF U308 ( .A(N605), .Y(N376) );
  INVX2TF U309 ( .A(N377), .Y(N603) );
  OR2X2TF U310 ( .A(N737), .B(STATE[3]), .Y(N1052) );
  NAND3X1TF U311 ( .A(STATE[2]), .B(N552), .C(STATE[1]), .Y(N737) );
  INVX2TF U312 ( .A(N1108), .Y(N1126) );
  AOI21X1TF U313 ( .A0(N672), .A1(N673), .B0(N671), .Y(N677) );
  AO21X1TF U314 ( .A0(N602), .A1(N1057), .B0(N787), .Y(N426) );
  OAI211XLTF U315 ( .A0(N728), .A1(N375), .B0(N733), .C0(N1130), .Y(
        NEXT_STATE[0]) );
  INVX2TF U316 ( .A(N264), .Y(N1131) );
  INVX2TF U317 ( .A(N1109), .Y(N1125) );
  INVX2TF U318 ( .A(N672), .Y(N674) );
  INVX2TF U319 ( .A(N673), .Y(N675) );
  NAND2X1TF U320 ( .A(N91), .B(N351), .Y(N684) );
  NAND2X1TF U321 ( .A(N351), .B(N335), .Y(N678) );
  NAND2X1TF U322 ( .A(N90), .B(N91), .Y(N689) );
  NAND2X1TF U323 ( .A(N90), .B(N335), .Y(N681) );
  OAI22X1TF U324 ( .A0(N671), .A1(N673), .B0(N672), .B1(N735), .Y(N653) );
  INVX2TF U325 ( .A(N651), .Y(N671) );
  INVX2TF U326 ( .A(N599), .Y(N1053) );
  INVX2TF U327 ( .A(N602), .Y(N1051) );
  OA21X2TF U328 ( .A0(N647), .A1(N393), .B0(N603), .Y(N602) );
  NAND2X1TF U329 ( .A(N356), .B(N360), .Y(N1032) );
  NOR2X4TF U330 ( .A(N1101), .B(N761), .Y(N1047) );
  NOR2BX2TF U331 ( .AN(CODE_TYPE[3]), .B(N2110), .Y(N611) );
  AND2X2TF U332 ( .A(N609), .B(N603), .Y(N599) );
  NOR2X2TF U333 ( .A(STATE[1]), .B(N733), .Y(N1133) );
  NAND3X1TF U334 ( .A(N307), .B(N1102), .C(N633), .Y(N1129) );
  INVX2TF U335 ( .A(N1104), .Y(N1130) );
  AOI21X2TF U336 ( .A0(N496), .A1(N268), .B0(N402), .Y(N600) );
  NOR2X1TF U337 ( .A(CODE_TYPE[3]), .B(N2110), .Y(N633) );
  AO22X1TF U338 ( .A0(N465), .A1(N601), .B0(N499), .B1(N268), .Y(N568) );
  AO22X1TF U339 ( .A0(N1062), .A1(CF), .B0(N589), .B1(CF_BUF), .Y(N4550) );
  OAI31XLTF U340 ( .A0(N348), .A1(STATE[3]), .A2(N552), .B0(N737), .Y(N729) );
  AO22X1TF U341 ( .A0(N264), .A1(N166), .B0(N1131), .B1(SMDR[11]), .Y(N4950)
         );
  AO22X1TF U342 ( .A0(N264), .A1(N177), .B0(N1131), .B1(SMDR[0]), .Y(N506) );
  AO22X1TF U343 ( .A0(N265), .A1(N176), .B0(N1131), .B1(SMDR[1]), .Y(N505) );
  AO22X1TF U344 ( .A0(N265), .A1(N170), .B0(N1131), .B1(SMDR[7]), .Y(N4990) );
  AO22X1TF U345 ( .A0(N264), .A1(N167), .B0(N1131), .B1(SMDR[10]), .Y(N4960)
         );
  AO22X1TF U346 ( .A0(N265), .A1(N162), .B0(N1131), .B1(SMDR[15]), .Y(N4910)
         );
  AO22X1TF U347 ( .A0(N265), .A1(N169), .B0(N1131), .B1(SMDR[8]), .Y(N4980) );
  AO22X1TF U348 ( .A0(N265), .A1(N164), .B0(N1131), .B1(SMDR[13]), .Y(N4930)
         );
  AO22X1TF U349 ( .A0(N265), .A1(N163), .B0(N1131), .B1(SMDR[14]), .Y(N4920)
         );
  AO22X1TF U350 ( .A0(N265), .A1(N165), .B0(N1131), .B1(SMDR[12]), .Y(N4940)
         );
  AO22X1TF U351 ( .A0(N264), .A1(N168), .B0(N1132), .B1(SMDR[9]), .Y(N4970) );
  AO22X1TF U352 ( .A0(N265), .A1(N175), .B0(N1132), .B1(SMDR[2]), .Y(N504) );
  AO22X1TF U353 ( .A0(N264), .A1(N173), .B0(N1132), .B1(SMDR[4]), .Y(N502) );
  AO22X1TF U354 ( .A0(N265), .A1(N171), .B0(N1132), .B1(SMDR[6]), .Y(N500) );
  AO22X1TF U355 ( .A0(N264), .A1(N172), .B0(N1132), .B1(SMDR[5]), .Y(N501) );
  AO22X1TF U356 ( .A0(N265), .A1(N174), .B0(N1132), .B1(SMDR[3]), .Y(N503) );
  AND4X1TF U357 ( .A(N633), .B(N1102), .C(N303), .D(N306), .Y(N158) );
  AOI22XLTF U358 ( .A0(N277), .A1(\IO_CONTROL[6] ), .B0(N2520), .B1(N32), .Y(
        N1245) );
  AOI22XLTF U359 ( .A0(N379), .A1(\IO_CONTROL[6] ), .B0(N2540), .B1(N32), .Y(
        N1173) );
  AOI22XLTF U360 ( .A0(N277), .A1(\IO_CONTROL[5] ), .B0(N2520), .B1(
        IO_DATAOUTB[5]), .Y(N1241) );
  AOI22XLTF U361 ( .A0(N379), .A1(\IO_CONTROL[5] ), .B0(N2540), .B1(
        IO_DATAOUTB[5]), .Y(N1169) );
  AOI22XLTF U362 ( .A0(N280), .A1(\IO_CONTROL[5] ), .B0(N256), .B1(
        IO_DATAOUTB[5]), .Y(N1313) );
  AOI22XLTF U363 ( .A0(N280), .A1(\IO_CONTROL[6] ), .B0(N256), .B1(N32), .Y(
        N1317) );
  INVX2TF U364 ( .A(N1092), .Y(N1085) );
  NAND2X1TF U365 ( .A(N1069), .B(N1104), .Y(N1075) );
  AND2X2TF U366 ( .A(N640), .B(N651), .Y(N719) );
  AOI221XLTF U367 ( .A0(N5670), .A1(NF), .B0(N634), .B1(N367), .C0(N346), .Y(
        N638) );
  INVX2TF U368 ( .A(N1139), .Y(N1138) );
  NAND2X2TF U369 ( .A(N1136), .B(N1135), .Y(N1139) );
  INVX2TF U370 ( .A(N1133), .Y(N1134) );
  NAND2BX1TF U371 ( .AN(N552), .B(N1135), .Y(N733) );
  INVX2TF U372 ( .A(N650), .Y(N735) );
  NOR2X2TF U373 ( .A(N5670), .B(N2000), .Y(N1102) );
  INVX2TF U374 ( .A(N632), .Y(N391) );
  INVX2TF U375 ( .A(N729), .Y(N734) );
  NOR2X1TF U376 ( .A(N723), .B(CPU_WAIT), .Y(N727) );
  OAI21X1TF U377 ( .A0(N332), .A1(N224), .B0(N1124), .Y(N4890) );
  AOI22X1TF U378 ( .A0(N382), .A1(\GR[5][1] ), .B0(N383), .B1(\GR[7][1] ), .Y(
        N1227) );
  AOI22X1TF U379 ( .A0(N380), .A1(\GR[5][1] ), .B0(N381), .B1(\GR[7][1] ), .Y(
        N1155) );
  OAI21X1TF U380 ( .A0(N334), .A1(N224), .B0(N1111), .Y(N476) );
  AOI22X1TF U381 ( .A0(N301), .A1(\GR[5][14] ), .B0(N1218), .B1(\GR[7][14] ), 
        .Y(N1279) );
  AOI22X1TF U382 ( .A0(N299), .A1(\GR[5][14] ), .B0(N1146), .B1(\GR[7][14] ), 
        .Y(N1207) );
  OAI21X1TF U383 ( .A0(N341), .A1(N224), .B0(N1117), .Y(N482) );
  AOI22X1TF U384 ( .A0(N301), .A1(\GR[5][8] ), .B0(N1218), .B1(\GR[7][8] ), 
        .Y(N1255) );
  AOI22X1TF U385 ( .A0(N299), .A1(\GR[5][8] ), .B0(N1146), .B1(\GR[7][8] ), 
        .Y(N1183) );
  OAI21X1TF U386 ( .A0(N349), .A1(N225), .B0(N1127), .Y(N4900) );
  AOI22X1TF U387 ( .A0(N382), .A1(\GR[5][0] ), .B0(N383), .B1(\GR[7][0] ), .Y(
        N1223) );
  AOI22X1TF U388 ( .A0(N380), .A1(\GR[5][0] ), .B0(N381), .B1(\GR[7][0] ), .Y(
        N1151) );
  OAI21X1TF U389 ( .A0(N342), .A1(N224), .B0(N1122), .Y(N4870) );
  AOI22X1TF U390 ( .A0(N382), .A1(\GR[5][3] ), .B0(N383), .B1(\GR[7][3] ), .Y(
        N1235) );
  AOI22X1TF U391 ( .A0(N380), .A1(\GR[5][3] ), .B0(N381), .B1(\GR[7][3] ), .Y(
        N1163) );
  OAI21X1TF U392 ( .A0(N338), .A1(N224), .B0(N1114), .Y(N479) );
  AOI22X1TF U393 ( .A0(N301), .A1(\GR[5][11] ), .B0(N383), .B1(\GR[7][11] ), 
        .Y(N1267) );
  AOI22X1TF U394 ( .A0(N299), .A1(\GR[5][11] ), .B0(N381), .B1(\GR[7][11] ), 
        .Y(N1195) );
  OAI21X1TF U395 ( .A0(N363), .A1(N224), .B0(N1119), .Y(N4840) );
  AOI22X1TF U396 ( .A0(N382), .A1(\GR[5][6] ), .B0(N383), .B1(\GR[7][6] ), .Y(
        N1247) );
  AOI22X1TF U397 ( .A0(N380), .A1(\GR[5][6] ), .B0(N381), .B1(\GR[7][6] ), .Y(
        N1175) );
  OAI21X1TF U398 ( .A0(N362), .A1(N224), .B0(N1121), .Y(N4860) );
  AOI22X1TF U399 ( .A0(N382), .A1(\GR[5][4] ), .B0(N383), .B1(\GR[7][4] ), .Y(
        N1239) );
  AOI22X1TF U400 ( .A0(N380), .A1(\GR[5][4] ), .B0(N381), .B1(\GR[7][4] ), .Y(
        N1167) );
  OAI21X1TF U401 ( .A0(N339), .A1(N224), .B0(N1123), .Y(N4880) );
  AOI22X1TF U402 ( .A0(N382), .A1(\GR[5][2] ), .B0(N383), .B1(\GR[7][2] ), .Y(
        N1231) );
  AOI22X1TF U403 ( .A0(N380), .A1(\GR[5][2] ), .B0(N381), .B1(\GR[7][2] ), .Y(
        N1159) );
  OAI21X1TF U404 ( .A0(N343), .A1(N225), .B0(N1118), .Y(N4830) );
  AOI22X1TF U405 ( .A0(N382), .A1(\GR[5][7] ), .B0(N383), .B1(\GR[7][7] ), .Y(
        N1251) );
  AOI22X1TF U406 ( .A0(N380), .A1(\GR[5][7] ), .B0(N381), .B1(\GR[7][7] ), .Y(
        N1179) );
  OAI21X1TF U407 ( .A0(N345), .A1(N225), .B0(N1112), .Y(N477) );
  AOI22X1TF U408 ( .A0(N301), .A1(\GR[5][13] ), .B0(N1218), .B1(\GR[7][13] ), 
        .Y(N1275) );
  AOI22X1TF U409 ( .A0(N299), .A1(\GR[5][13] ), .B0(N1146), .B1(\GR[7][13] ), 
        .Y(N1203) );
  OAI21X1TF U410 ( .A0(N333), .A1(N225), .B0(N1113), .Y(N478) );
  AOI22X1TF U411 ( .A0(N301), .A1(\GR[5][12] ), .B0(N1218), .B1(\GR[7][12] ), 
        .Y(N1271) );
  AOI22X1TF U413 ( .A0(N299), .A1(\GR[5][12] ), .B0(N1146), .B1(\GR[7][12] ), 
        .Y(N1199) );
  OAI21X1TF U414 ( .A0(N340), .A1(N225), .B0(N1116), .Y(N481) );
  AOI22X1TF U415 ( .A0(N382), .A1(\GR[5][9] ), .B0(N383), .B1(\GR[7][9] ), .Y(
        N1259) );
  AOI22X1TF U416 ( .A0(N380), .A1(\GR[5][9] ), .B0(N381), .B1(\GR[7][9] ), .Y(
        N1187) );
  OAI21X1TF U417 ( .A0(N350), .A1(N225), .B0(N1110), .Y(N475) );
  AOI22X1TF U418 ( .A0(N301), .A1(\GR[5][15] ), .B0(N1218), .B1(\GR[7][15] ), 
        .Y(N1283) );
  AOI22X1TF U419 ( .A0(N299), .A1(\GR[5][15] ), .B0(N1146), .B1(\GR[7][15] ), 
        .Y(N1211) );
  OAI21X1TF U420 ( .A0(N344), .A1(N225), .B0(N1115), .Y(N480) );
  AOI22X1TF U421 ( .A0(N301), .A1(\GR[5][10] ), .B0(N1218), .B1(\GR[7][10] ), 
        .Y(N1263) );
  AOI22X1TF U422 ( .A0(N299), .A1(\GR[5][10] ), .B0(N1146), .B1(\GR[7][10] ), 
        .Y(N1191) );
  OAI21X1TF U423 ( .A0(N361), .A1(N225), .B0(N1120), .Y(N4850) );
  AOI22X1TF U424 ( .A0(N382), .A1(\GR[5][5] ), .B0(N383), .B1(\GR[7][5] ), .Y(
        N1243) );
  AND3X2TF U425 ( .A(N94), .B(N92), .C(N93), .Y(N1218) );
  NOR3X1TF U426 ( .A(N93), .B(N371), .C(N337), .Y(N1217) );
  NOR3X4TF U427 ( .A(N92), .B(N93), .C(N337), .Y(N1215) );
  AOI22X1TF U428 ( .A0(N380), .A1(\GR[5][5] ), .B0(N381), .B1(\GR[7][5] ), .Y(
        N1171) );
  AND3X2TF U429 ( .A(N91), .B(N89), .C(N90), .Y(N1146) );
  NOR3X4TF U430 ( .A(N89), .B(N90), .C(N335), .Y(N1143) );
  OAI21X1TF U431 ( .A0(N1106), .A1(N1105), .B0(N1104), .Y(N1109) );
  OAI22X1TF U432 ( .A0(N1097), .A1(N1107), .B0(N1096), .B1(N1095), .Y(N1098)
         );
  INVX2TF U433 ( .A(N589), .Y(N1062) );
  OAI21X1TF U434 ( .A0(N352), .A1(N1094), .B0(N1091), .Y(N473) );
  AOI22X1TF U435 ( .A0(N384), .A1(\GR[5][1] ), .B0(N385), .B1(\GR[7][1] ), .Y(
        N1299) );
  OAI21X1TF U436 ( .A0(N370), .A1(N1094), .B0(N1093), .Y(N474) );
  AOI22X1TF U437 ( .A0(N384), .A1(\GR[5][0] ), .B0(N385), .B1(\GR[7][0] ), .Y(
        N1295) );
  OAI21X1TF U438 ( .A0(N336), .A1(N1094), .B0(N1090), .Y(N472) );
  AOI22X1TF U439 ( .A0(N384), .A1(\GR[5][2] ), .B0(N385), .B1(\GR[7][2] ), .Y(
        N1303) );
  OAI21X1TF U440 ( .A0(N259), .A1(N1094), .B0(N1089), .Y(N471) );
  AOI22X1TF U441 ( .A0(N384), .A1(\GR[5][3] ), .B0(N385), .B1(\GR[7][3] ), .Y(
        N1307) );
  OAI21X1TF U442 ( .A0(N259), .A1(N1075), .B0(N1074), .Y(N4630) );
  AOI22X1TF U443 ( .A0(N300), .A1(\GR[5][11] ), .B0(N1290), .B1(\GR[7][11] ), 
        .Y(N1339) );
  OAI21X1TF U444 ( .A0(N1075), .A1(N337), .B0(N1071), .Y(N4600) );
  AOI22X1TF U445 ( .A0(N300), .A1(\GR[5][14] ), .B0(N1290), .B1(\GR[7][14] ), 
        .Y(N1351) );
  OAI21X1TF U446 ( .A0(N577), .A1(N1085), .B0(N1076), .Y(N4640) );
  AOI22X1TF U447 ( .A0(N384), .A1(\GR[5][10] ), .B0(N1290), .B1(\GR[7][10] ), 
        .Y(N1335) );
  OAI21X1TF U448 ( .A0(N578), .A1(N1085), .B0(N1077), .Y(N4650) );
  AOI22X1TF U449 ( .A0(N384), .A1(\GR[5][9] ), .B0(N385), .B1(\GR[7][9] ), .Y(
        N1331) );
  OAI21X1TF U450 ( .A0(N582), .A1(N1085), .B0(N1082), .Y(N469) );
  AOI22X1TF U451 ( .A0(N300), .A1(\GR[5][5] ), .B0(N385), .B1(\GR[7][5] ), .Y(
        N1315) );
  OAI21X1TF U452 ( .A0(N583), .A1(N1085), .B0(N1084), .Y(N470) );
  AOI22X1TF U453 ( .A0(N300), .A1(\GR[5][4] ), .B0(N385), .B1(\GR[7][4] ), .Y(
        N1311) );
  OAI21X1TF U454 ( .A0(N575), .A1(N1085), .B0(N1073), .Y(N4620) );
  AOI22X1TF U455 ( .A0(N384), .A1(\GR[5][12] ), .B0(N1290), .B1(\GR[7][12] ), 
        .Y(N1343) );
  OAI21X1TF U456 ( .A0(N574), .A1(N1085), .B0(N1072), .Y(N4610) );
  AOI22X1TF U457 ( .A0(N384), .A1(\GR[5][13] ), .B0(N1290), .B1(\GR[7][13] ), 
        .Y(N1347) );
  OAI21X1TF U458 ( .A0(N581), .A1(N1085), .B0(N1081), .Y(N468) );
  AOI22X1TF U459 ( .A0(N300), .A1(\GR[5][6] ), .B0(N385), .B1(\GR[7][6] ), .Y(
        N1319) );
  OAI21X1TF U460 ( .A0(N580), .A1(N1085), .B0(N1080), .Y(N467) );
  NOR2X1TF U461 ( .A(N1086), .B(N1130), .Y(N1083) );
  AOI22X1TF U462 ( .A0(N300), .A1(\GR[5][7] ), .B0(N385), .B1(\GR[7][7] ), .Y(
        N1323) );
  OAI21X1TF U463 ( .A0(N579), .A1(N1085), .B0(N1079), .Y(N466) );
  AOI22X1TF U464 ( .A0(N384), .A1(\GR[5][8] ), .B0(N385), .B1(\GR[7][8] ), .Y(
        N1327) );
  INVX2TF U465 ( .A(N1075), .Y(N1078) );
  OAI21X1TF U466 ( .A0(N260), .A1(N1075), .B0(N1070), .Y(N4590) );
  OAI31X4TF U467 ( .A0(N1069), .A1(N1068), .A2(N1067), .B0(N1104), .Y(N1092)
         );
  AOI32X1TF U468 ( .A0(N1066), .A1(N1086), .A2(N1065), .B0(N29), .B1(N1086), 
        .Y(N1067) );
  AOI21X1TF U469 ( .A0(N359), .A1(N1103), .B0(N29), .Y(N1068) );
  AOI22X1TF U470 ( .A0(N300), .A1(\GR[5][15] ), .B0(N1290), .B1(\GR[7][15] ), 
        .Y(N1355) );
  AND3X2TF U471 ( .A(N97), .B(N95), .C(N96), .Y(N1290) );
  NOR3X1TF U472 ( .A(N96), .B(N370), .C(N336), .Y(N1289) );
  NOR3X4TF U473 ( .A(N95), .B(N96), .C(N336), .Y(N1287) );
  AOI21X1TF U474 ( .A0(N1095), .A1(N1054), .B0(N1096), .Y(N1069) );
  AOI211X1TF U475 ( .A0(N719), .A1(D_ADDR[8]), .B0(N718), .C0(N716), .Y(N717)
         );
  AOI211X1TF U476 ( .A0(N715), .A1(N366), .B0(N714), .C0(N713), .Y(N716) );
  NOR2X1TF U477 ( .A(N366), .B(N712), .Y(N718) );
  AOI211X1TF U478 ( .A0(N719), .A1(D_ADDR[6]), .B0(N708), .C0(N707), .Y(N722)
         );
  AOI211X1TF U479 ( .A0(N706), .A1(N365), .B0(N710), .C0(N713), .Y(N707) );
  NOR2X1TF U480 ( .A(N365), .B(N712), .Y(N708) );
  AOI211X1TF U481 ( .A0(N719), .A1(D_ADDR[4]), .B0(N702), .C0(N701), .Y(N724)
         );
  AOI211X1TF U482 ( .A0(N700), .A1(N364), .B0(N703), .C0(N713), .Y(N701) );
  NOR2X1TF U483 ( .A(N364), .B(N712), .Y(N702) );
  AOI22X1TF U484 ( .A0(N704), .A1(N709), .B0(I_ADDR[5]), .B1(N711), .Y(N705)
         );
  AOI21X1TF U485 ( .A0(I_ADDR[1]), .A1(N711), .B0(N641), .Y(N777) );
  INVX2TF U486 ( .A(N709), .Y(N713) );
  OAI32X1TF U487 ( .A0(N642), .A1(N714), .A2(I_ADDR[9]), .B0(N709), .B1(N642), 
        .Y(N776) );
  INVX2TF U488 ( .A(N712), .Y(N711) );
  OAI21X1TF U489 ( .A0(STATE[1]), .A1(N731), .B0(N639), .Y(N712) );
  OAI21X1TF U490 ( .A0(N640), .A1(N736), .B0(N651), .Y(N639) );
  NOR2X1TF U491 ( .A(N715), .B(N366), .Y(N714) );
  NOR2X1TF U492 ( .A(N706), .B(N365), .Y(N710) );
  NOR2X1TF U493 ( .A(N700), .B(N364), .Y(N703) );
  OAI32X1TF U494 ( .A0(N1107), .A1(N307), .A2(N638), .B0(N637), .B1(N1107), 
        .Y(N640) );
  AOI221X1TF U495 ( .A0(N636), .A1(ZF), .B0(N1102), .B1(N368), .C0(N635), .Y(
        N637) );
  INVX2TF U496 ( .A(N607), .Y(N1107) );
  AOI22X1TF U497 ( .A0(N1133), .A1(N1137), .B0(N259), .B1(N1134), .Y(N511) );
  INVX2TF U498 ( .A(I_DATAIN[3]), .Y(N1137) );
  OAI32X1TF U499 ( .A0(N606), .A1(N1104), .A2(N526), .B0(N730), .B1(N606), .Y(
        N961) );
  NOR2X1TF U500 ( .A(N737), .B(N1129), .Y(N595) );
  AOI2BB2X2TF U501 ( .B0(D_DATAIN[5]), .B1(N674), .A0N(N279), .A1N(N673), .Y(
        N695) );
  AOI22X2TF U502 ( .A0(REG_C[10]), .A1(N675), .B0(N674), .B1(D_DATAIN[2]), .Y(
        N692) );
  AOI22X2TF U503 ( .A0(REG_C[9]), .A1(N675), .B0(N674), .B1(D_DATAIN[1]), .Y(
        N691) );
  AOI22X2TF U504 ( .A0(REG_C[12]), .A1(N675), .B0(N674), .B1(D_DATAIN[4]), .Y(
        N694) );
  AOI22X2TF U505 ( .A0(REG_C[15]), .A1(N675), .B0(N674), .B1(D_DATAIN[7]), .Y(
        N697) );
  AOI22X2TF U506 ( .A0(REG_C[11]), .A1(N675), .B0(N674), .B1(D_DATAIN[3]), .Y(
        N693) );
  AOI22X2TF U507 ( .A0(REG_C[14]), .A1(N675), .B0(N674), .B1(D_DATAIN[6]), .Y(
        N696) );
  AOI22X2TF U508 ( .A0(D_ADDR[1]), .A1(N651), .B0(N650), .B1(D_DATAIN[0]), .Y(
        N662) );
  AOI22X2TF U509 ( .A0(N651), .A1(D_ADDR[3]), .B0(N650), .B1(D_DATAIN[2]), .Y(
        N664) );
  AOI22X2TF U510 ( .A0(N651), .A1(D_ADDR[5]), .B0(N650), .B1(D_DATAIN[4]), .Y(
        N666) );
  AOI22X2TF U511 ( .A0(N651), .A1(D_ADDR[7]), .B0(N650), .B1(D_DATAIN[6]), .Y(
        N668) );
  AOI22X2TF U512 ( .A0(N651), .A1(D_ADDR[4]), .B0(N650), .B1(D_DATAIN[3]), .Y(
        N665) );
  AOI22X2TF U513 ( .A0(D_ADDR[9]), .A1(N675), .B0(N674), .B1(D_DATAIN[0]), .Y(
        N690) );
  AOI22X2TF U514 ( .A0(N651), .A1(D_ADDR[2]), .B0(N650), .B1(D_DATAIN[1]), .Y(
        N663) );
  AOI22X2TF U515 ( .A0(N303), .A1(D_ADDR[8]), .B0(N650), .B1(D_DATAIN[7]), .Y(
        N669) );
  AOI22X2TF U516 ( .A0(N303), .A1(D_ADDR[6]), .B0(N650), .B1(D_DATAIN[5]), .Y(
        N667) );
  OAI211X1TF U517 ( .A0(N648), .A1(N1096), .B0(N647), .C0(N646), .Y(N649) );
  INVX2TF U518 ( .A(N610), .Y(N1096) );
  OAI211X1TF U519 ( .A0(N590), .A1(N1051), .B0(N1024), .C0(N1023), .Y(N446) );
  AOI22X1TF U520 ( .A0(IO_DATAINB[11]), .A1(N293), .B0(N599), .B1(N1060), .Y(
        N1023) );
  AOI22X1TF U521 ( .A0(IO_DATAINA[11]), .A1(N597), .B0(REG_C[11]), .B1(N1052), 
        .Y(N1024) );
  OAI211X1TF U522 ( .A0(N592), .A1(N1051), .B0(N981), .C0(N980), .Y(N438) );
  AOI22X1TF U523 ( .A0(IO_DATAINA[7]), .A1(N217), .B0(N599), .B1(N1061), .Y(
        N980) );
  AOI22X1TF U524 ( .A0(IO_DATAINB[7]), .A1(N293), .B0(D_ADDR[8]), .B1(N1052), 
        .Y(N981) );
  INVX2TF U525 ( .A(N586), .Y(N585) );
  OAI211X1TF U526 ( .A0(N593), .A1(N1053), .B0(N977), .C0(N976), .Y(N436) );
  AOI22X1TF U527 ( .A0(IO_DATAINA[6]), .A1(N217), .B0(N602), .B1(N1061), .Y(
        N976) );
  AOI21X1TF U528 ( .A0(N376), .A1(N970), .B0(N581), .Y(N975) );
  AOI22X1TF U529 ( .A0(REG_A[6]), .A1(N608), .B0(N387), .B1(N363), .Y(N970) );
  AOI21X1TF U530 ( .A0(N386), .A1(N581), .B0(N1047), .Y(N4490) );
  AOI22X1TF U531 ( .A0(IO_DATAINB[6]), .A1(N293), .B0(D_ADDR[7]), .B1(N377), 
        .Y(N977) );
  OAI211X1TF U532 ( .A0(N593), .A1(N1051), .B0(N966), .C0(N965), .Y(N434) );
  AOI22X1TF U533 ( .A0(IO_DATAINA[5]), .A1(N217), .B0(N599), .B1(N1059), .Y(
        N965) );
  AOI22X1TF U534 ( .A0(IO_DATAINB[5]), .A1(N293), .B0(D_ADDR[6]), .B1(N1052), 
        .Y(N966) );
  AOI211X1TF U535 ( .A0(N488), .A1(N268), .B0(N447), .C0(N964), .Y(N593) );
  OAI22X1TF U536 ( .A0(N830), .A1(N361), .B0(N829), .B1(N994), .Y(N964) );
  AOI21X1TF U537 ( .A0(N388), .A1(N582), .B0(N1047), .Y(N830) );
  INVX2TF U538 ( .A(N445), .Y(N447) );
  AOI211X1TF U539 ( .A0(N828), .A1(N443), .B0(N963), .C0(N441), .Y(N445) );
  AOI211X1TF U540 ( .A0(N386), .A1(N361), .B0(N437), .C0(N1044), .Y(N439) );
  NOR2X1TF U541 ( .A(N1013), .B(N361), .Y(N437) );
  OAI22X1TF U542 ( .A0(N991), .A1(N979), .B0(N995), .B1(N992), .Y(N963) );
  OAI211X1TF U543 ( .A0(N590), .A1(N1053), .B0(N1027), .C0(N1026), .Y(N448) );
  AOI22X1TF U544 ( .A0(IO_DATAINB[12]), .A1(N293), .B0(N602), .B1(N1025), .Y(
        N1026) );
  INVX2TF U545 ( .A(N598), .Y(N1025) );
  AOI22X1TF U546 ( .A0(IO_DATAINA[12]), .A1(N217), .B0(REG_C[12]), .B1(N377), 
        .Y(N1027) );
  AOI21X1TF U547 ( .A0(N494), .A1(N268), .B0(N539), .Y(N590) );
  OAI211X1TF U548 ( .A0(N553), .A1(N1021), .B0(N1020), .C0(N537), .Y(N538) );
  AOI21X1TF U549 ( .A0(N1018), .A1(N1019), .B0(N1022), .Y(N537) );
  OAI32X1TF U550 ( .A0(N338), .A1(N357), .A2(REG_B[11]), .B0(N614), .B1(N338), 
        .Y(N1022) );
  OAI22X1TF U551 ( .A0(N1017), .A1(N1032), .B0(N1016), .B1(N1015), .Y(N1018)
         );
  OAI21X1TF U552 ( .A0(N1014), .A1(N1044), .B0(REG_B[11]), .Y(N1020) );
  AOI22X1TF U553 ( .A0(REG_A[11]), .A1(N1013), .B0(N357), .B1(N338), .Y(N1014)
         );
  OAI21X1TF U554 ( .A0(N588), .A1(N1051), .B0(N587), .Y(N4540) );
  AOI22X1TF U555 ( .A0(N586), .A1(N599), .B0(REG_C[15]), .B1(N377), .Y(N587)
         );
  AOI21X1TF U556 ( .A0(N463), .A1(N546), .B0(N541), .Y(N542) );
  OAI211X1TF U557 ( .A0(N1050), .A1(N553), .B0(N1049), .C0(N540), .Y(N541) );
  AOI32X1TF U558 ( .A0(N387), .A1(REG_A[14]), .A2(N573), .B0(N1047), .B1(
        REG_A[14]), .Y(N1048) );
  AOI22X1TF U559 ( .A0(REG_A[14]), .A1(N608), .B0(N387), .B1(N334), .Y(N1029)
         );
  AOI22X1TF U560 ( .A0(N1046), .A1(N1045), .B0(N1044), .B1(REG_B[14]), .Y(
        N1049) );
  NOR2X1TF U561 ( .A(N972), .B(N971), .Y(N1045) );
  AOI211X1TF U562 ( .A0(N1043), .A1(N1042), .B0(N1041), .C0(N1040), .Y(N1050)
         );
  OAI22X1TF U563 ( .A0(N1039), .A1(N1038), .B0(N1037), .B1(N1036), .Y(N1040)
         );
  AOI31X1TF U564 ( .A0(N1035), .A1(N1034), .A2(N1033), .B0(N1032), .Y(N1041)
         );
  AOI22X1TF U565 ( .A0(N302), .A1(REG_A[14]), .B0(N1030), .B1(REG_A[12]), .Y(
        N1035) );
  OAI211X1TF U566 ( .A0(N591), .A1(N1051), .B0(N1008), .C0(N1007), .Y(N444) );
  AOI22X1TF U567 ( .A0(IO_DATAINB[10]), .A1(N293), .B0(N599), .B1(N1056), .Y(
        N1007) );
  AOI22X1TF U568 ( .A0(IO_DATAINA[10]), .A1(N217), .B0(REG_C[10]), .B1(N377), 
        .Y(N1008) );
  OAI211X1TF U569 ( .A0(N594), .A1(N1053), .B0(N786), .C0(N785), .Y(N787) );
  AOI22X1TF U570 ( .A0(N293), .A1(IO_DATAINB[1]), .B0(N5950), .B1(IO_STATUS[1]), .Y(N785) );
  AOI22X1TF U571 ( .A0(IO_DATAINA[1]), .A1(N217), .B0(D_ADDR[2]), .B1(N377), 
        .Y(N786) );
  AOI21X1TF U572 ( .A0(IO_DATAINA[0]), .A1(N597), .B0(N563), .Y(N564) );
  OAI211X1TF U573 ( .A0(N594), .A1(N1051), .B0(N562), .C0(N561), .Y(N563) );
  AOI22X1TF U574 ( .A0(N596), .A1(IO_DATAINB[0]), .B0(D_ADDR[1]), .B1(N377), 
        .Y(N562) );
  AOI21X1TF U575 ( .A0(N421), .A1(REG_A[0]), .B0(N420), .Y(N594) );
  OAI211X1TF U576 ( .A0(N972), .A1(N746), .B0(N745), .C0(N419), .Y(N420) );
  AOI21X1TF U577 ( .A0(N449), .A1(N378), .B0(N418), .Y(N419) );
  OAI211X1TF U578 ( .A0(REG_A[0]), .A1(N357), .B0(N416), .C0(N376), .Y(N417)
         );
  OAI31X1TF U579 ( .A0(N744), .A1(N743), .A2(N758), .B0(N988), .Y(N745) );
  NOR2X1TF U580 ( .A(N339), .B(N30), .Y(N743) );
  NOR2X1TF U581 ( .A(N332), .B(N756), .Y(N744) );
  OAI21X1TF U582 ( .A0(N198), .A1(N357), .B0(N544), .Y(N421) );
  INVX2TF U583 ( .A(N591), .Y(N1060) );
  AND2X2TF U584 ( .A(N536), .B(N535), .Y(N591) );
  AOI21X1TF U585 ( .A0(N459), .A1(N378), .B0(N534), .Y(N535) );
  AOI21X1TF U586 ( .A0(N1042), .A1(N612), .B0(N531), .Y(N532) );
  OAI22X1TF U587 ( .A0(N530), .A1(N577), .B0(N755), .B1(N344), .Y(N531) );
  AOI21X1TF U588 ( .A0(N388), .A1(N577), .B0(N1047), .Y(N755) );
  OAI22X1TF U589 ( .A0(N1039), .A1(N983), .B0(N1037), .B1(N973), .Y(N760) );
  NOR2X1TF U590 ( .A(N2090), .B(N342), .Y(N758) );
  AND2X2TF U591 ( .A(N412), .B(N411), .Y(N598) );
  AOI21X1TF U592 ( .A0(N461), .A1(N378), .B0(N410), .Y(N411) );
  NOR2X1TF U593 ( .A(N791), .B(N741), .Y(N403) );
  AOI221X1TF U594 ( .A0(N386), .A1(N333), .B0(N608), .B1(REG_A[12]), .C0(N1044), .Y(N630) );
  OAI211X1TF U595 ( .A0(N994), .A1(N991), .B0(N401), .C0(N625), .Y(N402) );
  AOI211X1TF U596 ( .A0(N604), .A1(N1000), .B0(N624), .C0(N623), .Y(N625) );
  OAI22X1TF U597 ( .A0(N574), .A1(N622), .B0(N621), .B1(N345), .Y(N623) );
  AOI21X1TF U598 ( .A0(N574), .A1(N388), .B0(N626), .Y(N621) );
  OAI21X1TF U599 ( .A0(N762), .A1(N968), .B0(N614), .Y(N626) );
  AOI221X1TF U600 ( .A0(N608), .A1(REG_A[13]), .B0(N387), .B1(N345), .C0(N1044), .Y(N622) );
  OAI22X1TF U601 ( .A0(N827), .A1(N620), .B0(N619), .B1(N968), .Y(N624) );
  AOI211X1TF U602 ( .A0(N1030), .A1(REG_A[11]), .B0(N814), .C0(N810), .Y(N619)
         );
  AOI22X1TF U603 ( .A0(REG_B[2]), .A1(N778), .B0(N996), .B1(N356), .Y(N827) );
  OAI22X1TF U604 ( .A0(N550), .A1(N572), .B0(N549), .B1(N968), .Y(N551) );
  AOI211X1TF U605 ( .A0(N1030), .A1(REG_A[13]), .B0(N548), .C0(N768), .Y(N549)
         );
  NOR2X1TF U606 ( .A(N756), .B(N334), .Y(N548) );
  AOI21X1TF U607 ( .A0(N608), .A1(REG_A[15]), .B0(N547), .Y(N550) );
  OAI21X1TF U608 ( .A0(N357), .A1(REG_A[15]), .B0(N376), .Y(N547) );
  AOI21X1TF U609 ( .A0(N386), .A1(N572), .B0(N545), .Y(N557) );
  INVX2TF U610 ( .A(N544), .Y(N545) );
  AOI21X1TF U611 ( .A0(N612), .A1(N302), .B0(N815), .Y(N544) );
  OAI211X1TF U612 ( .A0(N592), .A1(N1053), .B0(N990), .C0(N989), .Y(N440) );
  AOI22X1TF U613 ( .A0(IO_DATAINA[8]), .A1(N217), .B0(N602), .B1(N1055), .Y(
        N989) );
  AOI22X1TF U614 ( .A0(IO_DATAINB[8]), .A1(N293), .B0(D_ADDR[9]), .B1(N377), 
        .Y(N990) );
  OAI211X1TF U615 ( .A0(N576), .A1(N1053), .B0(N571), .C0(N570), .Y(N584) );
  OR2X2TF U616 ( .A(N826), .B(N435), .Y(N1059) );
  AOI21X1TF U617 ( .A0(N831), .A1(N987), .B0(N427), .Y(N433) );
  AOI21X1TF U618 ( .A0(N386), .A1(N583), .B0(N1047), .Y(N423) );
  OAI22X1TF U619 ( .A0(N986), .A1(N979), .B0(N973), .B1(N982), .Y(N825) );
  AOI21X1TF U620 ( .A0(N376), .A1(N823), .B0(N583), .Y(N826) );
  AOI22X1TF U621 ( .A0(REG_A[4]), .A1(N608), .B0(N387), .B1(N362), .Y(N823) );
  AOI22X1TF U622 ( .A0(N596), .A1(IO_DATAINB[4]), .B0(D_ADDR[5]), .B1(N1052), 
        .Y(N571) );
  OAI211X1TF U623 ( .A0(N576), .A1(N1051), .B0(N5680), .C0(N566), .Y(N569) );
  AOI22X1TF U624 ( .A0(N596), .A1(IO_DATAINB[3]), .B0(D_ADDR[4]), .B1(N377), 
        .Y(N5680) );
  OAI211X1TF U625 ( .A0(N2120), .A1(N361), .B0(N806), .C0(N805), .Y(N807) );
  OAI211X1TF U626 ( .A0(N1017), .A1(N979), .B0(N820), .C0(N819), .Y(N821) );
  AOI221X1TF U627 ( .A0(N342), .A1(N387), .B0(REG_A[3]), .B1(N608), .C0(N816), 
        .Y(N817) );
  OAI31X1TF U628 ( .A0(N356), .A1(N972), .A2(N1015), .B0(N376), .Y(N816) );
  AOI22X1TF U629 ( .A0(N831), .A1(N978), .B0(N486), .B1(N267), .Y(N820) );
  NOR2X1TF U630 ( .A(N2100), .B(N344), .Y(N814) );
  AOI211X1TF U631 ( .A0(N302), .A1(REG_A[11]), .B0(N810), .C0(N809), .Y(N1017)
         );
  OAI22X1TF U632 ( .A0(N345), .A1(N30), .B0(N2100), .B1(N334), .Y(N809) );
  NOR2X1TF U633 ( .A(N756), .B(N333), .Y(N810) );
  OAI211X1TF U634 ( .A0(N2100), .A1(N349), .B0(N748), .C0(N773), .Y(N1010) );
  AOI22X1TF U635 ( .A0(N1031), .A1(REG_A[3]), .B0(REG_A[1]), .B1(N2130), .Y(
        N748) );
  OAI211X1TF U636 ( .A0(N1006), .A1(N1051), .B0(N1005), .C0(N1004), .Y(N442)
         );
  AOI22X1TF U637 ( .A0(IO_DATAINA[9]), .A1(N597), .B0(N599), .B1(N1055), .Y(
        N1004) );
  OAI211X1TF U638 ( .A0(N2100), .A1(N332), .B0(N628), .C0(N792), .Y(N984) );
  AOI22X1TF U639 ( .A0(N1031), .A1(REG_A[4]), .B0(REG_A[2]), .B1(N2130), .Y(
        N628) );
  INVX2TF U640 ( .A(N742), .Y(N986) );
  OAI211X1TF U641 ( .A0(N333), .A1(N762), .B0(N1033), .C0(N627), .Y(N742) );
  AOI22X1TF U642 ( .A0(N808), .A1(REG_A[15]), .B0(N2130), .B1(REG_A[14]), .Y(
        N627) );
  INVX2TF U643 ( .A(N824), .Y(N982) );
  NOR2X1TF U644 ( .A(N762), .B(N349), .Y(N824) );
  INVX2TF U645 ( .A(N357), .Y(N388) );
  NOR2X1TF U646 ( .A(N30), .B(N344), .Y(N741) );
  INVX2TF U647 ( .A(N994), .Y(N988) );
  AOI22X1TF U648 ( .A0(IO_DATAINB[9]), .A1(N293), .B0(REG_C[9]), .B1(N1052), 
        .Y(N1005) );
  INVX2TF U649 ( .A(N1056), .Y(N1006) );
  OAI211X1TF U650 ( .A0(N578), .A1(N1003), .B0(N1002), .C0(N1001), .Y(N1056)
         );
  AOI211X1TF U651 ( .A0(N612), .A1(N1000), .B0(N999), .C0(N998), .Y(N1001) );
  OAI211X1TF U652 ( .A0(N973), .A1(N528), .B0(N527), .C0(N525), .Y(N998) );
  OAI211X1TF U653 ( .A0(N2100), .A1(N339), .B0(N618), .C0(N806), .Y(N996) );
  AOI22X1TF U654 ( .A0(N1031), .A1(REG_A[5]), .B0(REG_A[3]), .B1(N2130), .Y(
        N618) );
  INVX2TF U655 ( .A(N604), .Y(N973) );
  AND2X2TF U656 ( .A(N613), .B(N1043), .Y(N604) );
  OAI22X1TF U657 ( .A0(N995), .A1(N994), .B0(N993), .B1(N340), .Y(N999) );
  AOI21X1TF U658 ( .A0(N387), .A1(N578), .B0(N1047), .Y(N993) );
  INVX2TF U659 ( .A(N831), .Y(N992) );
  AOI221X1TF U660 ( .A0(N386), .A1(N340), .B0(N292), .B1(REG_A[9]), .C0(N1044), 
        .Y(N1003) );
  AOI22X1TF U661 ( .A0(N599), .A1(N1057), .B0(N602), .B1(N1058), .Y(N802) );
  AOI22X1TF U662 ( .A0(N378), .A1(N451), .B0(N485), .B1(N267), .Y(N422) );
  AOI211X1TF U663 ( .A0(N831), .A1(N969), .B0(N800), .C0(N799), .Y(N801) );
  OAI22X1TF U664 ( .A0(N798), .A1(N339), .B0(N797), .B1(N356), .Y(N799) );
  AOI221X1TF U665 ( .A0(N386), .A1(N339), .B0(N608), .B1(REG_A[2]), .C0(N1044), 
        .Y(N797) );
  INVX2TF U666 ( .A(N1013), .Y(N608) );
  INVX2TF U667 ( .A(N357), .Y(N386) );
  AOI21X1TF U668 ( .A0(N387), .A1(N356), .B0(N815), .Y(N798) );
  OAI22X1TF U669 ( .A0(N796), .A1(N994), .B0(N360), .B1(N795), .Y(N800) );
  AOI211X1TF U670 ( .A0(REG_A[10]), .A1(N302), .B0(N750), .C0(N749), .Y(N967)
         );
  OAI22X1TF U671 ( .A0(N345), .A1(N2090), .B0(N30), .B1(N333), .Y(N749) );
  NOR2X1TF U672 ( .A(N756), .B(N338), .Y(N750) );
  AOI211X1TF U673 ( .A0(REG_A[4]), .A1(N1030), .B0(N794), .C0(N793), .Y(N796)
         );
  NOR2X1TF U674 ( .A(N2090), .B(N361), .Y(N793) );
  INVX2TF U675 ( .A(N792), .Y(N794) );
  NOR2X1TF U676 ( .A(N2100), .B(N340), .Y(N791) );
  NOR2X1TF U677 ( .A(N1016), .B(N972), .Y(N831) );
  OR2X2TF U678 ( .A(N1032), .B(N553), .Y(N968) );
  INVX2TF U679 ( .A(N613), .Y(N553) );
  AOI21X1TF U680 ( .A0(N1031), .A1(REG_A[2]), .B0(N757), .Y(N1039) );
  OAI22X1TF U681 ( .A0(N349), .A1(N30), .B0(N332), .B1(N756), .Y(N757) );
  AND2X2TF U682 ( .A(N5670), .B(N358), .Y(N393) );
  OAI211X1TF U683 ( .A0(N784), .A1(N972), .B0(N783), .C0(N782), .Y(N1057) );
  AOI32X1TF U684 ( .A0(N387), .A1(REG_A[1]), .A2(N355), .B0(N815), .B1(
        REG_A[1]), .Y(N782) );
  OAI21X1TF U685 ( .A0(N762), .A1(N994), .B0(N614), .Y(N815) );
  INVX2TF U686 ( .A(N1047), .Y(N614) );
  INVX2TF U687 ( .A(N357), .Y(N387) );
  AOI211X1TF U688 ( .A0(REG_B[1]), .A1(N781), .B0(N780), .C0(N779), .Y(N783)
         );
  AOI22X1TF U689 ( .A0(N413), .A1(N443), .B0(N484), .B1(N267), .Y(N414) );
  INVX2TF U690 ( .A(N1054), .Y(N394) );
  AND2X2TF U691 ( .A(N613), .B(N360), .Y(N443) );
  NOR2X2TF U692 ( .A(CODE_TYPE[1]), .B(N389), .Y(N613) );
  INVX2TF U693 ( .A(N1088), .Y(N389) );
  INVX2TF U694 ( .A(N997), .Y(N413) );
  AOI221X1TF U695 ( .A0(N198), .A1(N349), .B0(N354), .B1(N332), .C0(REG_B[1]), 
        .Y(N778) );
  OR2X2TF U696 ( .A(N400), .B(N399), .Y(N546) );
  AND2X2TF U697 ( .A(N611), .B(N1097), .Y(N601) );
  NOR2X1TF U698 ( .A(N2000), .B(CODE_TYPE[1]), .Y(N1097) );
  NOR2X1TF U699 ( .A(N397), .B(N1100), .Y(N400) );
  NOR2X1TF U700 ( .A(N358), .B(N648), .Y(N1100) );
  NOR2X1TF U701 ( .A(N634), .B(N2000), .Y(N636) );
  AOI31X1TF U702 ( .A0(N775), .A1(N774), .A2(N773), .B0(N994), .Y(N780) );
  NAND2X2TF U703 ( .A(N1046), .B(N1019), .Y(N994) );
  INVX2TF U704 ( .A(N972), .Y(N1019) );
  INVX2TF U705 ( .A(N1032), .Y(N1046) );
  INVX2TF U706 ( .A(N756), .Y(N747) );
  INVX2TF U707 ( .A(N30), .Y(N1030) );
  AOI21X1TF U708 ( .A0(N607), .A1(N392), .B0(N391), .Y(N605) );
  INVX2TF U709 ( .A(N1095), .Y(N392) );
  AND2X2TF U710 ( .A(CODE_TYPE[3]), .B(N29), .Y(N607) );
  OR2X2TF U711 ( .A(N1064), .B(N1101), .Y(N1013) );
  INVX2TF U712 ( .A(N611), .Y(N1101) );
  NOR2X2TF U713 ( .A(N346), .B(N648), .Y(N1063) );
  INVX2TF U714 ( .A(N772), .Y(N784) );
  INVX2TF U715 ( .A(N1009), .Y(N1036) );
  NOR2X2TF U716 ( .A(REG_B[2]), .B(N360), .Y(N1009) );
  NOR4X1TF U717 ( .A(N771), .B(N770), .C(N769), .D(N768), .Y(N995) );
  NOR2X1TF U718 ( .A(N333), .B(N2090), .Y(N768) );
  NOR2X1TF U719 ( .A(N756), .B(N344), .Y(N769) );
  NOR2X1TF U720 ( .A(N30), .B(N338), .Y(N770) );
  NOR2X1TF U721 ( .A(N762), .B(N340), .Y(N771) );
  INVX2TF U722 ( .A(N767), .Y(N1038) );
  NOR2X1TF U723 ( .A(N356), .B(N360), .Y(N767) );
  AOI21X1TF U724 ( .A0(REG_A[13]), .A1(N302), .B0(N616), .Y(N991) );
  OAI22X1TF U725 ( .A0(N30), .A1(N350), .B0(N756), .B1(N334), .Y(N616) );
  INVX2TF U726 ( .A(N1043), .Y(N1016) );
  NOR4X1TF U727 ( .A(N766), .B(N765), .C(N764), .D(N763), .Y(N829) );
  NOR2X1TF U728 ( .A(N2100), .B(N341), .Y(N763) );
  NOR2X1TF U729 ( .A(N756), .B(N363), .Y(N764) );
  NOR2X1TF U730 ( .A(N30), .B(N343), .Y(N765) );
  NOR2X1TF U731 ( .A(N762), .B(N361), .Y(N766) );
  INVX2TF U732 ( .A(N1031), .Y(N762) );
  INVX2TF U733 ( .A(N633), .Y(N390) );
  AOI22X1TF U734 ( .A0(N293), .A1(IO_DATAINB[2]), .B0(N5950), .B1(IO_STATUS[2]), .Y(N803) );
  NOR2X1TF U735 ( .A(N415), .B(N761), .Y(N5950) );
  INVX2TF U736 ( .A(N1103), .Y(N615) );
  AOI22X1TF U737 ( .A0(IO_DATAINA[2]), .A1(N597), .B0(D_ADDR[3]), .B1(N377), 
        .Y(N804) );
  NOR3X4TF U738 ( .A(N415), .B(N1103), .C(CODE_TYPE[1]), .Y(N597) );
  AOI22X1TF U739 ( .A0(N277), .A1(\IO_CONTROL[1] ), .B0(N2520), .B1(
        IO_DATAOUTB[1]), .Y(N1225) );
  AOI22X1TF U740 ( .A0(N298), .A1(\IO_CONTROL[1] ), .B0(N255), .B1(
        IO_DATAOUTB[1]), .Y(N1153) );
  AOI22X1TF U741 ( .A0(N282), .A1(\GR[0][1] ), .B0(N258), .B1(N33), .Y(N1152)
         );
  AOI22X1TF U742 ( .A0(N278), .A1(N1357), .B0(N2530), .B1(N1368), .Y(N1277) );
  AOI22X1TF U743 ( .A0(N227), .A1(\GR[0][14] ), .B0(N275), .B1(N1365), .Y(
        N1276) );
  AOI22X1TF U744 ( .A0(N298), .A1(N1357), .B0(N255), .B1(N1368), .Y(N1205) );
  AOI22X1TF U745 ( .A0(N282), .A1(\GR[0][14] ), .B0(N261), .B1(N1365), .Y(
        N1204) );
  AOI22X1TF U746 ( .A0(N277), .A1(N1363), .B0(N2520), .B1(IO_DATAOUTB[8]), .Y(
        N1253) );
  AOI22X1TF U747 ( .A0(N298), .A1(N1363), .B0(N255), .B1(IO_DATAOUTB[8]), .Y(
        N1181) );
  AOI22X1TF U748 ( .A0(N282), .A1(\GR[0][8] ), .B0(N258), .B1(N40), .Y(N1180)
         );
  AOI22X1TF U749 ( .A0(N277), .A1(\IO_CONTROL[0] ), .B0(N2520), .B1(
        IO_DATAOUTB[0]), .Y(N1221) );
  AOI22X1TF U750 ( .A0(N1143), .A1(IO_OFFSET[0]), .B0(N269), .B1(\GR[6][0] ), 
        .Y(N1150) );
  AOI22X1TF U751 ( .A0(N379), .A1(\IO_CONTROL[0] ), .B0(N2540), .B1(
        IO_DATAOUTB[0]), .Y(N1149) );
  AOI22X1TF U752 ( .A0(N282), .A1(\GR[0][0] ), .B0(N258), .B1(IO_DATAOUTA[0]), 
        .Y(N1148) );
  AOI22X1TF U753 ( .A0(N278), .A1(\IO_CONTROL[3] ), .B0(N2520), .B1(N38), .Y(
        N1233) );
  AOI22X1TF U754 ( .A0(N226), .A1(\GR[0][3] ), .B0(N275), .B1(IO_DATAOUTA[3]), 
        .Y(N1232) );
  AOI22X1TF U755 ( .A0(N379), .A1(\IO_CONTROL[3] ), .B0(N2540), .B1(N38), .Y(
        N1161) );
  AOI22X1TF U756 ( .A0(N283), .A1(\GR[0][3] ), .B0(N258), .B1(IO_DATAOUTA[3]), 
        .Y(N1160) );
  AOI22X1TF U757 ( .A0(N277), .A1(N1360), .B0(N2520), .B1(N44), .Y(N1265) );
  AOI22X1TF U758 ( .A0(N227), .A1(\GR[0][11] ), .B0(N276), .B1(IO_DATAOUTA[11]), .Y(N1264) );
  AOI22X1TF U759 ( .A0(N379), .A1(N1360), .B0(N2540), .B1(N44), .Y(N1193) );
  AOI22X1TF U760 ( .A0(N283), .A1(\GR[0][11] ), .B0(N258), .B1(IO_DATAOUTA[11]), .Y(N1192) );
  AOI22X1TF U761 ( .A0(N1215), .A1(IO_OFFSET[6]), .B0(N273), .B1(\GR[6][6] ), 
        .Y(N1246) );
  AOI22X1TF U762 ( .A0(N282), .A1(\GR[0][6] ), .B0(N258), .B1(N36), .Y(N1172)
         );
  AOI22X1TF U763 ( .A0(N310), .A1(IO_OFFSET[4]), .B0(N274), .B1(\GR[6][4] ), 
        .Y(N1238) );
  AOI22X1TF U764 ( .A0(N278), .A1(\IO_CONTROL[4] ), .B0(N2530), .B1(N39), .Y(
        N1237) );
  AOI22X1TF U765 ( .A0(N227), .A1(\GR[0][4] ), .B0(N276), .B1(N35), .Y(N1236)
         );
  AOI22X1TF U766 ( .A0(N1143), .A1(IO_OFFSET[4]), .B0(N270), .B1(\GR[6][4] ), 
        .Y(N1166) );
  AOI22X1TF U767 ( .A0(N379), .A1(\IO_CONTROL[4] ), .B0(N2540), .B1(N39), .Y(
        N1165) );
  AOI22X1TF U768 ( .A0(N283), .A1(\GR[0][4] ), .B0(N261), .B1(N35), .Y(N1164)
         );
  AOI22X1TF U769 ( .A0(N310), .A1(IO_OFFSET[2]), .B0(N273), .B1(\GR[6][2] ), 
        .Y(N1230) );
  AOI22X1TF U770 ( .A0(N1143), .A1(IO_OFFSET[2]), .B0(N269), .B1(\GR[6][2] ), 
        .Y(N1158) );
  AOI22X1TF U771 ( .A0(N310), .A1(IO_OFFSET[7]), .B0(N274), .B1(\GR[6][7] ), 
        .Y(N1250) );
  AOI22X1TF U772 ( .A0(N278), .A1(\IO_CONTROL[7] ), .B0(N2530), .B1(
        IO_DATAOUTB[7]), .Y(N1249) );
  AOI22X1TF U773 ( .A0(N227), .A1(\GR[0][7] ), .B0(N276), .B1(N37), .Y(N1248)
         );
  AOI22X1TF U774 ( .A0(N308), .A1(IO_OFFSET[7]), .B0(N270), .B1(\GR[6][7] ), 
        .Y(N1178) );
  AOI22X1TF U775 ( .A0(N379), .A1(\IO_CONTROL[7] ), .B0(N2540), .B1(
        IO_DATAOUTB[7]), .Y(N1177) );
  AOI22X1TF U776 ( .A0(N283), .A1(\GR[0][7] ), .B0(N261), .B1(N37), .Y(N1176)
         );
  AOI22X1TF U777 ( .A0(N310), .A1(N1372), .B0(N274), .B1(\GR[6][13] ), .Y(
        N1274) );
  AOI22X1TF U778 ( .A0(N278), .A1(N1358), .B0(N2530), .B1(N1369), .Y(N1273) );
  AOI22X1TF U779 ( .A0(N227), .A1(\GR[0][13] ), .B0(N276), .B1(N1366), .Y(
        N1272) );
  AOI22X1TF U780 ( .A0(N308), .A1(N1372), .B0(N270), .B1(\GR[6][13] ), .Y(
        N1202) );
  AOI22X1TF U781 ( .A0(N298), .A1(N1358), .B0(N255), .B1(N1369), .Y(N1201) );
  AOI22X1TF U782 ( .A0(N283), .A1(\GR[0][13] ), .B0(N261), .B1(N1366), .Y(
        N1200) );
  AOI22X1TF U783 ( .A0(N310), .A1(N1373), .B0(N274), .B1(\GR[6][12] ), .Y(
        N1270) );
  AOI22X1TF U784 ( .A0(N278), .A1(N1359), .B0(N2530), .B1(IO_DATAOUTB[12]), 
        .Y(N1269) );
  AOI22X1TF U785 ( .A0(N227), .A1(\GR[0][12] ), .B0(N276), .B1(N43), .Y(N1268)
         );
  AOI22X1TF U786 ( .A0(N308), .A1(N1373), .B0(N270), .B1(\GR[6][12] ), .Y(
        N1198) );
  AOI22X1TF U787 ( .A0(N298), .A1(N1359), .B0(N255), .B1(IO_DATAOUTB[12]), .Y(
        N1197) );
  AOI22X1TF U788 ( .A0(N283), .A1(\GR[0][12] ), .B0(N261), .B1(N43), .Y(N1196)
         );
  AOI22X1TF U789 ( .A0(N1215), .A1(IO_OFFSET[9]), .B0(N274), .B1(\GR[6][9] ), 
        .Y(N1258) );
  AOI22X1TF U790 ( .A0(N278), .A1(N1362), .B0(N2530), .B1(IO_DATAOUTB[9]), .Y(
        N1257) );
  AOI22X1TF U791 ( .A0(N227), .A1(\GR[0][9] ), .B0(N276), .B1(N41), .Y(N1256)
         );
  AOI22X1TF U792 ( .A0(N308), .A1(IO_OFFSET[9]), .B0(N270), .B1(\GR[6][9] ), 
        .Y(N1186) );
  AOI22X1TF U793 ( .A0(N379), .A1(N1362), .B0(N255), .B1(IO_DATAOUTB[9]), .Y(
        N1185) );
  AOI22X1TF U794 ( .A0(N283), .A1(\GR[0][9] ), .B0(N261), .B1(N41), .Y(N1184)
         );
  AOI22X1TF U795 ( .A0(N310), .A1(N1370), .B0(N274), .B1(\GR[6][15] ), .Y(
        N1282) );
  AOI22X1TF U796 ( .A0(N278), .A1(N1356), .B0(N2530), .B1(N1367), .Y(N1281) );
  AOI22X1TF U797 ( .A0(N227), .A1(\GR[0][15] ), .B0(N276), .B1(N1364), .Y(
        N1280) );
  AOI22X1TF U798 ( .A0(N308), .A1(N1370), .B0(N270), .B1(\GR[6][15] ), .Y(
        N1210) );
  AOI22X1TF U799 ( .A0(N298), .A1(N1356), .B0(N255), .B1(N1367), .Y(N1209) );
  AOI22X1TF U800 ( .A0(N283), .A1(\GR[0][15] ), .B0(N261), .B1(N1364), .Y(
        N1208) );
  AOI22X1TF U801 ( .A0(N310), .A1(N1375), .B0(N274), .B1(\GR[6][10] ), .Y(
        N1262) );
  AOI22X1TF U802 ( .A0(N278), .A1(N1361), .B0(N2530), .B1(IO_DATAOUTB[10]), 
        .Y(N1261) );
  AOI22X1TF U803 ( .A0(N227), .A1(\GR[0][10] ), .B0(N276), .B1(N42), .Y(N1260)
         );
  AOI22X1TF U804 ( .A0(N308), .A1(N1375), .B0(N270), .B1(\GR[6][10] ), .Y(
        N1190) );
  AOI22X1TF U805 ( .A0(N298), .A1(N1361), .B0(N255), .B1(IO_DATAOUTB[10]), .Y(
        N1189) );
  AOI22X1TF U806 ( .A0(N283), .A1(\GR[0][10] ), .B0(N261), .B1(N42), .Y(N1188)
         );
  AOI22X1TF U807 ( .A0(N1215), .A1(IO_OFFSET[5]), .B0(N274), .B1(\GR[6][5] ), 
        .Y(N1242) );
  AOI22X1TF U808 ( .A0(N308), .A1(IO_OFFSET[5]), .B0(N270), .B1(\GR[6][5] ), 
        .Y(N1170) );
  AOI22X1TF U809 ( .A0(N282), .A1(\GR[0][5] ), .B0(N258), .B1(IO_DATAOUTA[5]), 
        .Y(N1168) );
  AOI22X1TF U810 ( .A0(REG_B[1]), .A1(N1092), .B0(N222), .B1(N253), .Y(N1091)
         );
  AOI22X1TF U811 ( .A0(N280), .A1(\IO_CONTROL[1] ), .B0(N256), .B1(
        IO_DATAOUTB[1]), .Y(N1297) );
  AOI22X1TF U812 ( .A0(N284), .A1(\GR[0][1] ), .B0(N262), .B1(N33), .Y(N1296)
         );
  AOI22X1TF U813 ( .A0(N198), .A1(N1092), .B0(N222), .B1(N254), .Y(N1093) );
  AOI22X1TF U814 ( .A0(N280), .A1(\IO_CONTROL[0] ), .B0(N256), .B1(
        IO_DATAOUTB[0]), .Y(N1293) );
  AOI22X1TF U815 ( .A0(N284), .A1(\GR[0][0] ), .B0(N262), .B1(IO_DATAOUTA[0]), 
        .Y(N1292) );
  AOI22X1TF U816 ( .A0(REG_B[2]), .A1(N1092), .B0(N222), .B1(N252), .Y(N1090)
         );
  AOI22X1TF U817 ( .A0(REG_B[3]), .A1(N1092), .B0(N222), .B1(N251), .Y(N1089)
         );
  AOI22X1TF U818 ( .A0(N280), .A1(\IO_CONTROL[3] ), .B0(N257), .B1(N38), .Y(
        N1305) );
  AOI22X1TF U819 ( .A0(N284), .A1(\GR[0][3] ), .B0(N263), .B1(IO_DATAOUTA[3]), 
        .Y(N1304) );
  AOI22X1TF U820 ( .A0(N243), .A1(N221), .B0(N1092), .B1(REG_B[11]), .Y(N1074)
         );
  AOI22X1TF U821 ( .A0(N309), .A1(N1374), .B0(N272), .B1(\GR[6][11] ), .Y(
        N1338) );
  AOI22X1TF U822 ( .A0(N281), .A1(N1360), .B0(N257), .B1(N44), .Y(N1337) );
  AOI22X1TF U823 ( .A0(N285), .A1(\GR[0][11] ), .B0(N263), .B1(IO_DATAOUTA[11]), .Y(N1336) );
  AOI22X1TF U824 ( .A0(N240), .A1(N221), .B0(N1092), .B1(REG_B[14]), .Y(N1071)
         );
  AOI22X1TF U825 ( .A0(N309), .A1(N1371), .B0(N272), .B1(\GR[6][14] ), .Y(
        N1350) );
  AOI22X1TF U826 ( .A0(N281), .A1(N1357), .B0(N257), .B1(N1368), .Y(N1349) );
  AOI22X1TF U827 ( .A0(N285), .A1(\GR[0][14] ), .B0(N263), .B1(N1365), .Y(
        N1348) );
  AOI22X1TF U828 ( .A0(N1078), .A1(N97), .B0(N222), .B1(N244), .Y(N1076) );
  AOI22X1TF U829 ( .A0(N1287), .A1(N1375), .B0(N272), .B1(\GR[6][10] ), .Y(
        N1334) );
  AOI22X1TF U830 ( .A0(N281), .A1(N1361), .B0(N257), .B1(IO_DATAOUTB[10]), .Y(
        N1333) );
  AOI22X1TF U831 ( .A0(N285), .A1(\GR[0][10] ), .B0(N262), .B1(N42), .Y(N1332)
         );
  AOI22X1TF U832 ( .A0(N1078), .A1(N96), .B0(N222), .B1(N245), .Y(N1077) );
  AOI22X1TF U833 ( .A0(N280), .A1(N1362), .B0(N256), .B1(IO_DATAOUTB[9]), .Y(
        N1329) );
  AOI22X1TF U834 ( .A0(N284), .A1(\GR[0][9] ), .B0(N262), .B1(N41), .Y(N1328)
         );
  AOI22X1TF U835 ( .A0(N221), .A1(N249), .B0(N93), .B1(N1083), .Y(N1082) );
  AOI22X1TF U836 ( .A0(N309), .A1(IO_OFFSET[5]), .B0(N272), .B1(\GR[6][5] ), 
        .Y(N1314) );
  AOI22X1TF U837 ( .A0(N285), .A1(\GR[0][5] ), .B0(N263), .B1(IO_DATAOUTA[5]), 
        .Y(N1312) );
  AOI22X1TF U838 ( .A0(N221), .A1(N250), .B0(N92), .B1(N1083), .Y(N1084) );
  AOI22X1TF U839 ( .A0(N309), .A1(IO_OFFSET[4]), .B0(N272), .B1(\GR[6][4] ), 
        .Y(N1310) );
  AOI22X1TF U840 ( .A0(N281), .A1(\IO_CONTROL[4] ), .B0(N257), .B1(N39), .Y(
        N1309) );
  AOI22X1TF U841 ( .A0(N285), .A1(\GR[0][4] ), .B0(N263), .B1(N35), .Y(N1308)
         );
  AOI22X1TF U842 ( .A0(N1078), .A1(N92), .B0(N221), .B1(N242), .Y(N1073) );
  AOI22X1TF U843 ( .A0(N280), .A1(N1359), .B0(N256), .B1(IO_DATAOUTB[12]), .Y(
        N1341) );
  AOI22X1TF U844 ( .A0(N284), .A1(\GR[0][12] ), .B0(N262), .B1(N43), .Y(N1340)
         );
  AOI22X1TF U845 ( .A0(N1078), .A1(N93), .B0(N221), .B1(N241), .Y(N1072) );
  AOI22X1TF U846 ( .A0(N1287), .A1(N1372), .B0(N271), .B1(\GR[6][13] ), .Y(
        N1346) );
  AOI22X1TF U847 ( .A0(N281), .A1(N1358), .B0(N256), .B1(N1369), .Y(N1345) );
  AOI22X1TF U848 ( .A0(N284), .A1(\GR[0][13] ), .B0(N262), .B1(N1366), .Y(
        N1344) );
  AOI22X1TF U849 ( .A0(N221), .A1(N248), .B0(N94), .B1(N1083), .Y(N1081) );
  AOI22X1TF U850 ( .A0(N309), .A1(IO_OFFSET[6]), .B0(N272), .B1(\GR[6][6] ), 
        .Y(N1318) );
  AOI22X1TF U851 ( .A0(N285), .A1(\GR[0][6] ), .B0(N263), .B1(N36), .Y(N1316)
         );
  AOI22X1TF U852 ( .A0(N247), .A1(N221), .B0(N1083), .B1(N372), .Y(N1080) );
  AOI22X1TF U853 ( .A0(N309), .A1(IO_OFFSET[7]), .B0(N272), .B1(\GR[6][7] ), 
        .Y(N1322) );
  AOI22X1TF U854 ( .A0(N281), .A1(\IO_CONTROL[7] ), .B0(N257), .B1(
        IO_DATAOUTB[7]), .Y(N1321) );
  AOI22X1TF U855 ( .A0(N285), .A1(\GR[0][7] ), .B0(N263), .B1(N37), .Y(N1320)
         );
  AOI22X1TF U856 ( .A0(N1078), .A1(N95), .B0(N222), .B1(N246), .Y(N1079) );
  AOI22X1TF U857 ( .A0(N1287), .A1(IO_OFFSET[8]), .B0(N271), .B1(\GR[6][8] ), 
        .Y(N1326) );
  AOI22X1TF U858 ( .A0(N281), .A1(N1363), .B0(N257), .B1(IO_DATAOUTB[8]), .Y(
        N1325) );
  AOI22X1TF U859 ( .A0(N284), .A1(\GR[0][8] ), .B0(N262), .B1(N40), .Y(N1324)
         );
  AOI22X1TF U860 ( .A0(N309), .A1(N1370), .B0(N272), .B1(\GR[6][15] ), .Y(
        N1354) );
  AOI22X1TF U861 ( .A0(N281), .A1(N1356), .B0(N257), .B1(N1367), .Y(N1353) );
  AOI22X1TF U862 ( .A0(N285), .A1(\GR[0][15] ), .B0(N263), .B1(N1364), .Y(
        N1352) );
  OAI32XLTF U863 ( .A0(STATE[3]), .A1(STATE[2]), .A2(START), .B0(N552), .B1(
        STATE[3]), .Y(N631) );
  AOI22XLTF U864 ( .A0(STATE[3]), .A1(STATE[2]), .B0(N1135), .B1(N727), .Y(
        N728) );
  NOR3XLTF U865 ( .A(N90), .B(N369), .C(N335), .Y(N1145) );
  NOR3XLTF U866 ( .A(N91), .B(N90), .C(N369), .Y(N1142) );
  MXI2X1TF U867 ( .A(N588), .B(N367), .S0(N1062), .Y(N4560) );
  AOI22XLTF U868 ( .A0(N1135), .A1(N552), .B0(N1136), .B1(N348), .Y(N643) );
  OAI222X1TF U869 ( .A0(N1053), .A1(N600), .B0(N374), .B1(N603), .C0(N1051), 
        .C1(N585), .Y(N4520) );
  NAND3BX1TF U870 ( .AN(N521), .B(N516), .C(N4580), .Y(N1061) );
  AOI2BB1X1TF U871 ( .A0N(N1037), .A1N(N968), .B0(N975), .Y(N4580) );
  NAND2X1TF U872 ( .A(N489), .B(N268), .Y(N516) );
  NAND3BX1TF U873 ( .AN(N974), .B(N4530), .C(N4510), .Y(N521) );
  AOI2BB2X1TF U874 ( .B0(N455), .B1(N378), .A0N(N992), .A1N(N967), .Y(N4510)
         );
  AOI2BB2X1TF U875 ( .B0(N969), .B1(N988), .A0N(N4490), .A1N(N363), .Y(N4530)
         );
  AO21X1TF U876 ( .A0(N460), .A1(N546), .B0(N538), .Y(N539) );
  OAI2BB1X1TF U877 ( .A0N(N268), .A1N(N497), .B0(N542), .Y(N586) );
  OA21XLTF U878 ( .A0(N573), .A1(N1029), .B0(N1048), .Y(N540) );
  NAND2X1TF U879 ( .A(IO_STATUS[0]), .B(N5950), .Y(N561) );
  AO22X1TF U880 ( .A0(N417), .A1(N198), .B0(N483), .B1(N267), .Y(N418) );
  NAND2X1TF U881 ( .A(N608), .B(REG_A[0]), .Y(N416) );
  NAND2BX1TF U882 ( .AN(N760), .B(N533), .Y(N534) );
  OA21XLTF U883 ( .A0(N795), .A1(REG_B[3]), .B0(N532), .Y(N533) );
  AOI2BB1X1TF U884 ( .A0N(N1013), .A1N(N344), .B0(N529), .Y(N530) );
  OAI2BB1X1TF U885 ( .A0N(N344), .A1N(N388), .B0(N376), .Y(N529) );
  NAND2X1TF U886 ( .A(N493), .B(N267), .Y(N536) );
  NAND3X1TF U887 ( .A(N409), .B(N408), .C(N407), .Y(N410) );
  NAND2X1TF U888 ( .A(N406), .B(REG_A[12]), .Y(N407) );
  AO21X1TF U889 ( .A0(N386), .A1(N575), .B0(N626), .Y(N406) );
  AOI2BB1X1TF U890 ( .A0N(N994), .A1N(N986), .B0(N405), .Y(N408) );
  NAND2BX1TF U891 ( .AN(N750), .B(N403), .Y(N404) );
  NAND2BX1TF U892 ( .AN(N629), .B(N613), .Y(N409) );
  NAND2X1TF U893 ( .A(N495), .B(N267), .Y(N412) );
  NAND2X1TF U894 ( .A(N462), .B(N546), .Y(N401) );
  AOI2BB1X1TF U895 ( .A0N(N554), .A1N(N553), .B0(N551), .Y(N555) );
  AOI222XLTF U896 ( .A0(N1010), .A1(N767), .B0(N1011), .B1(N1009), .C0(N1012), 
        .C1(N1043), .Y(N554) );
  NAND2X1TF U897 ( .A(N1059), .B(N602), .Y(N570) );
  NAND4BX1TF U898 ( .AN(N825), .B(N433), .C(N431), .D(N429), .Y(N435) );
  NAND2X1TF U899 ( .A(N984), .B(N612), .Y(N429) );
  NAND2X1TF U900 ( .A(N487), .B(N267), .Y(N431) );
  OAI2BB1X1TF U901 ( .A0N(N988), .A1N(N822), .B0(N425), .Y(N427) );
  AOI2BB2X1TF U902 ( .B0(N378), .B1(N453), .A0N(N423), .A1N(N362), .Y(N425) );
  NAND2X1TF U903 ( .A(N1058), .B(N599), .Y(N566) );
  AO22X1TF U904 ( .A0(N546), .A1(N452), .B0(N807), .B1(N988), .Y(N543) );
  NAND3BX1TF U905 ( .AN(N997), .B(N613), .C(REG_B[3]), .Y(N525) );
  NAND2X1TF U906 ( .A(N458), .B(N378), .Y(N527) );
  OAI2BB1X1TF U907 ( .A0N(N450), .A1N(N378), .B0(N414), .Y(N779) );
  NAND2X1TF U908 ( .A(N610), .B(N394), .Y(N395) );
  NAND2X1TF U909 ( .A(CODE_TYPE[1]), .B(N1102), .Y(N1054) );
  MXI2X1TF U910 ( .A(N1103), .B(N2000), .S0(CODE_TYPE[1]), .Y(N396) );
  NAND2BX1TF U911 ( .AN(N601), .B(N398), .Y(N399) );
  NAND2X1TF U912 ( .A(N607), .B(CODE_TYPE[1]), .Y(N398) );
  OA21XLTF U913 ( .A0(N636), .A1(N358), .B0(N617), .Y(N397) );
  ADDHXLTF U914 ( .A(REG_A[0]), .B(REG_B[0]), .CO(ADD_X_300_3_N22), .S(N449)
         );
  CLKBUFX2TF U915 ( .A(N1218), .Y(N383) );
  CLKBUFX2TF U916 ( .A(N1146), .Y(N381) );
  CLKBUFX2TF U917 ( .A(N1290), .Y(N385) );
  OAI2BB1X1TF U918 ( .A0N(N2000), .A1N(N648), .B0(N359), .Y(N617) );
  NAND2X1TF U919 ( .A(N808), .B(REG_A[6]), .Y(N805) );
  NAND2X1TF U920 ( .A(N747), .B(REG_A[8]), .Y(N813) );
  NAND4BBX1TF U921 ( .AN(N771), .BN(N765), .C(N805), .D(N813), .Y(N1000) );
  NAND2X1TF U922 ( .A(REG_A[4]), .B(N747), .Y(N806) );
  NAND2X1TF U923 ( .A(N613), .B(REG_B[3]), .Y(N620) );
  NAND3X1TF U924 ( .A(N5670), .B(N346), .C(N306), .Y(N1095) );
  NAND2X1TF U925 ( .A(REG_A[13]), .B(N747), .Y(N1033) );
  NAND2X1TF U926 ( .A(N1031), .B(REG_A[8]), .Y(N740) );
  NAND2X1TF U927 ( .A(N2130), .B(REG_A[6]), .Y(N738) );
  NAND2X1TF U928 ( .A(N747), .B(REG_A[7]), .Y(N790) );
  NAND4BX1TF U929 ( .AN(N793), .B(N740), .C(N738), .D(N790), .Y(N985) );
  NAND2X1TF U930 ( .A(REG_A[3]), .B(N747), .Y(N792) );
  AOI222XLTF U931 ( .A0(N985), .A1(N1043), .B0(N824), .B1(N767), .C0(N984), 
        .C1(N1009), .Y(N629) );
  OAI222X1TF U932 ( .A0(N1051), .A1(N600), .B0(N1053), .B1(N598), .C0(N279), 
        .C1(N603), .Y(N4500) );
  NAND3X1TF U933 ( .A(I_ADDR[2]), .B(I_ADDR[1]), .C(I_ADDR[3]), .Y(N700) );
  NAND2X1TF U934 ( .A(I_ADDR[5]), .B(N703), .Y(N706) );
  NAND2X1TF U935 ( .A(N710), .B(I_ADDR[7]), .Y(N715) );
  NAND3X1TF U936 ( .A(N651), .B(N714), .C(I_ADDR[9]), .Y(N736) );
  AO22X1TF U937 ( .A0(I_ADDR[0]), .A1(SMDR[8]), .B0(N347), .B1(SMDR[0]), .Y(
        D_DATAOUT[0]) );
  AO22X1TF U938 ( .A0(I_ADDR[0]), .A1(SMDR[9]), .B0(N347), .B1(SMDR[1]), .Y(
        D_DATAOUT[1]) );
  AO22X1TF U939 ( .A0(I_ADDR[0]), .A1(SMDR[10]), .B0(N347), .B1(SMDR[2]), .Y(
        D_DATAOUT[2]) );
  AO22X1TF U940 ( .A0(I_ADDR[0]), .A1(SMDR[11]), .B0(N347), .B1(SMDR[3]), .Y(
        D_DATAOUT[3]) );
  AO22X1TF U941 ( .A0(I_ADDR[0]), .A1(SMDR[12]), .B0(N347), .B1(SMDR[4]), .Y(
        D_DATAOUT[4]) );
  AO22X1TF U942 ( .A0(I_ADDR[0]), .A1(SMDR[13]), .B0(N347), .B1(SMDR[5]), .Y(
        D_DATAOUT[5]) );
  AO22X1TF U943 ( .A0(I_ADDR[0]), .A1(SMDR[14]), .B0(N347), .B1(SMDR[6]), .Y(
        D_DATAOUT[6]) );
  AO22X1TF U944 ( .A0(I_ADDR[0]), .A1(SMDR[15]), .B0(N347), .B1(SMDR[7]), .Y(
        D_DATAOUT[7]) );
  NAND3X1TF U945 ( .A(N552), .B(N1135), .C(START), .Y(N731) );
  AOI2BB2X1TF U946 ( .B0(CF), .B1(N761), .A0N(N1063), .A1N(CF), .Y(N635) );
  OAI2BB2XLTF U947 ( .B0(I_ADDR[1]), .B1(N713), .A0N(D_ADDR[1]), .A1N(N719), 
        .Y(N641) );
  AO22X1TF U948 ( .A0(I_ADDR[9]), .A1(N711), .B0(N719), .B1(D_ADDR[9]), .Y(
        N642) );
  NAND2X1TF U949 ( .A(N552), .B(STATE[1]), .Y(N645) );
  NAND2BX1TF U950 ( .AN(N645), .B(N1135), .Y(N730) );
  OAI221XLTF U951 ( .A0(N307), .A1(N610), .B0(N306), .B1(N358), .C0(N5670), 
        .Y(N646) );
  AOI2BB2X1TF U952 ( .B0(N2470), .B1(N662), .A0N(\GR[0][0] ), .A1N(N2460), .Y(
        N960) );
  AOI2BB2X1TF U953 ( .B0(N2470), .B1(N663), .A0N(\GR[0][1] ), .A1N(N2460), .Y(
        N959) );
  AOI2BB2X1TF U954 ( .B0(N2470), .B1(N664), .A0N(\GR[0][2] ), .A1N(N2460), .Y(
        N958) );
  AOI2BB2X1TF U955 ( .B0(N2470), .B1(N665), .A0N(\GR[0][3] ), .A1N(N2460), .Y(
        N957) );
  AOI2BB2X1TF U956 ( .B0(N2470), .B1(N666), .A0N(\GR[0][4] ), .A1N(N2460), .Y(
        N956) );
  AOI2BB2X1TF U957 ( .B0(N2470), .B1(N667), .A0N(\GR[0][5] ), .A1N(N2460), .Y(
        N955) );
  AOI2BB2X1TF U958 ( .B0(N2470), .B1(N668), .A0N(\GR[0][6] ), .A1N(N2460), .Y(
        N954) );
  AOI2BB2X1TF U959 ( .B0(N2470), .B1(N669), .A0N(\GR[0][7] ), .A1N(N2460), .Y(
        N953) );
  AOI2BB2X1TF U960 ( .B0(N296), .B1(N662), .A0N(\IO_CONTROL[0] ), .A1N(N654), 
        .Y(N952) );
  AOI2BB2X1TF U961 ( .B0(N296), .B1(N663), .A0N(\IO_CONTROL[1] ), .A1N(N654), 
        .Y(N951) );
  AOI2BB2X1TF U962 ( .B0(N296), .B1(N664), .A0N(\IO_CONTROL[2] ), .A1N(N654), 
        .Y(N950) );
  AOI2BB2X1TF U963 ( .B0(N296), .B1(N665), .A0N(\IO_CONTROL[3] ), .A1N(N654), 
        .Y(N949) );
  AOI2BB2X1TF U964 ( .B0(N296), .B1(N666), .A0N(\IO_CONTROL[4] ), .A1N(N654), 
        .Y(N948) );
  AOI2BB2X1TF U965 ( .B0(N296), .B1(N667), .A0N(\IO_CONTROL[5] ), .A1N(N654), 
        .Y(N947) );
  AOI2BB2X1TF U966 ( .B0(N296), .B1(N668), .A0N(\IO_CONTROL[6] ), .A1N(N654), 
        .Y(N946) );
  AOI2BB2X1TF U967 ( .B0(N296), .B1(N669), .A0N(\IO_CONTROL[7] ), .A1N(N654), 
        .Y(N945) );
  AOI2BB2X1TF U968 ( .B0(N297), .B1(N662), .A0N(IO_DATAOUTA[0]), .A1N(N655), 
        .Y(N944) );
  AOI2BB2X1TF U969 ( .B0(N297), .B1(N663), .A0N(N33), .A1N(N655), .Y(N943) );
  AOI2BB2X1TF U970 ( .B0(N297), .B1(N664), .A0N(N34), .A1N(N655), .Y(N942) );
  AOI2BB2X1TF U971 ( .B0(N297), .B1(N665), .A0N(IO_DATAOUTA[3]), .A1N(N655), 
        .Y(N941) );
  AOI2BB2X1TF U972 ( .B0(N297), .B1(N666), .A0N(N35), .A1N(N655), .Y(N940) );
  AOI2BB2X1TF U973 ( .B0(N297), .B1(N667), .A0N(IO_DATAOUTA[5]), .A1N(N655), 
        .Y(N939) );
  AOI2BB2X1TF U974 ( .B0(N297), .B1(N668), .A0N(N36), .A1N(N655), .Y(N938) );
  AOI2BB2X1TF U975 ( .B0(N297), .B1(N669), .A0N(N37), .A1N(N655), .Y(N937) );
  AOI2BB2X1TF U976 ( .B0(N2430), .B1(N662), .A0N(IO_DATAOUTB[0]), .A1N(N2420), 
        .Y(N936) );
  AOI2BB2X1TF U977 ( .B0(N2430), .B1(N663), .A0N(IO_DATAOUTB[1]), .A1N(N2420), 
        .Y(N935) );
  AOI2BB2X1TF U978 ( .B0(N2430), .B1(N664), .A0N(IO_DATAOUTB[2]), .A1N(N2420), 
        .Y(N934) );
  AOI2BB2X1TF U979 ( .B0(N2430), .B1(N665), .A0N(N38), .A1N(N2420), .Y(N933)
         );
  AOI2BB2X1TF U980 ( .B0(N2430), .B1(N666), .A0N(N39), .A1N(N2420), .Y(N932)
         );
  AOI2BB2X1TF U981 ( .B0(N2430), .B1(N667), .A0N(IO_DATAOUTB[5]), .A1N(N2420), 
        .Y(N931) );
  AOI2BB2X1TF U982 ( .B0(N2430), .B1(N668), .A0N(N32), .A1N(N2420), .Y(N930)
         );
  AOI2BB2X1TF U983 ( .B0(N2430), .B1(N669), .A0N(IO_DATAOUTB[7]), .A1N(N2420), 
        .Y(N929) );
  AOI2BB2X1TF U984 ( .B0(N2410), .B1(N662), .A0N(IO_OFFSET[0]), .A1N(N2400), 
        .Y(N928) );
  AOI2BB2X1TF U985 ( .B0(N2410), .B1(N663), .A0N(IO_OFFSET[1]), .A1N(N2400), 
        .Y(N927) );
  AOI2BB2X1TF U986 ( .B0(N2410), .B1(N664), .A0N(IO_OFFSET[2]), .A1N(N2400), 
        .Y(N926) );
  AOI2BB2X1TF U987 ( .B0(N2410), .B1(N665), .A0N(IO_OFFSET[3]), .A1N(N2400), 
        .Y(N925) );
  AOI2BB2X1TF U988 ( .B0(N2410), .B1(N666), .A0N(IO_OFFSET[4]), .A1N(N2400), 
        .Y(N924) );
  AOI2BB2X1TF U989 ( .B0(N2410), .B1(N667), .A0N(IO_OFFSET[5]), .A1N(N2400), 
        .Y(N923) );
  AOI2BB2X1TF U990 ( .B0(N2410), .B1(N668), .A0N(IO_OFFSET[6]), .A1N(N2400), 
        .Y(N922) );
  AOI2BB2X1TF U991 ( .B0(N2410), .B1(N669), .A0N(IO_OFFSET[7]), .A1N(N2400), 
        .Y(N921) );
  AOI2BB2X1TF U992 ( .B0(N2490), .B1(N662), .A0N(\GR[5][0] ), .A1N(N2480), .Y(
        N920) );
  AOI2BB2X1TF U993 ( .B0(N2490), .B1(N663), .A0N(\GR[5][1] ), .A1N(N2480), .Y(
        N919) );
  AOI2BB2X1TF U994 ( .B0(N2490), .B1(N664), .A0N(\GR[5][2] ), .A1N(N2480), .Y(
        N918) );
  AOI2BB2X1TF U995 ( .B0(N2490), .B1(N665), .A0N(\GR[5][3] ), .A1N(N2480), .Y(
        N917) );
  AOI2BB2X1TF U996 ( .B0(N2490), .B1(N666), .A0N(\GR[5][4] ), .A1N(N2480), .Y(
        N916) );
  AOI2BB2X1TF U997 ( .B0(N2490), .B1(N667), .A0N(\GR[5][5] ), .A1N(N2480), .Y(
        N915) );
  AOI2BB2X1TF U998 ( .B0(N2490), .B1(N668), .A0N(\GR[5][6] ), .A1N(N2480), .Y(
        N914) );
  AOI2BB2X1TF U999 ( .B0(N2490), .B1(N669), .A0N(\GR[5][7] ), .A1N(N2480), .Y(
        N913) );
  AOI2BB2X1TF U1000 ( .B0(N2510), .B1(N662), .A0N(\GR[6][0] ), .A1N(N2500), 
        .Y(N912) );
  AOI2BB2X1TF U1001 ( .B0(N2510), .B1(N663), .A0N(\GR[6][1] ), .A1N(N2500), 
        .Y(N911) );
  AOI2BB2X1TF U1002 ( .B0(N2510), .B1(N664), .A0N(\GR[6][2] ), .A1N(N2500), 
        .Y(N910) );
  AOI2BB2X1TF U1003 ( .B0(N2510), .B1(N665), .A0N(\GR[6][3] ), .A1N(N2500), 
        .Y(N909) );
  AOI2BB2X1TF U1004 ( .B0(N2510), .B1(N666), .A0N(\GR[6][4] ), .A1N(N2500), 
        .Y(N908) );
  AOI2BB2X1TF U1005 ( .B0(N2510), .B1(N667), .A0N(\GR[6][5] ), .A1N(N2500), 
        .Y(N907) );
  AOI2BB2X1TF U1006 ( .B0(N2510), .B1(N668), .A0N(\GR[6][6] ), .A1N(N2500), 
        .Y(N906) );
  AOI2BB2X1TF U1007 ( .B0(N2510), .B1(N669), .A0N(\GR[6][7] ), .A1N(N2500), 
        .Y(N905) );
  AOI2BB2X1TF U1008 ( .B0(N2450), .B1(N662), .A0N(\GR[7][0] ), .A1N(N2440), 
        .Y(N904) );
  AOI2BB2X1TF U1009 ( .B0(N2450), .B1(N663), .A0N(\GR[7][1] ), .A1N(N2440), 
        .Y(N903) );
  AOI2BB2X1TF U1010 ( .B0(N2450), .B1(N664), .A0N(\GR[7][2] ), .A1N(N2440), 
        .Y(N902) );
  AOI2BB2X1TF U1011 ( .B0(N2450), .B1(N665), .A0N(\GR[7][3] ), .A1N(N2440), 
        .Y(N901) );
  AOI2BB2X1TF U1012 ( .B0(N2450), .B1(N666), .A0N(\GR[7][4] ), .A1N(N2440), 
        .Y(N900) );
  AOI2BB2X1TF U1013 ( .B0(N2450), .B1(N667), .A0N(\GR[7][5] ), .A1N(N2440), 
        .Y(N899) );
  AOI2BB2X1TF U1014 ( .B0(N2450), .B1(N668), .A0N(\GR[7][6] ), .A1N(N2440), 
        .Y(N898) );
  AOI2BB2X1TF U1015 ( .B0(N2450), .B1(N669), .A0N(\GR[7][7] ), .A1N(N2440), 
        .Y(N897) );
  AOI2BB2X1TF U1016 ( .B0(N2390), .B1(N690), .A0N(\GR[0][8] ), .A1N(N238), .Y(
        N896) );
  AOI2BB2X1TF U1017 ( .B0(N2390), .B1(N691), .A0N(\GR[0][9] ), .A1N(N238), .Y(
        N895) );
  AOI2BB2X1TF U1018 ( .B0(N2390), .B1(N692), .A0N(\GR[0][10] ), .A1N(N238), 
        .Y(N894) );
  AOI2BB2X1TF U1019 ( .B0(N2390), .B1(N693), .A0N(\GR[0][11] ), .A1N(N238), 
        .Y(N893) );
  AOI2BB2X1TF U1020 ( .B0(N2390), .B1(N694), .A0N(\GR[0][12] ), .A1N(N238), 
        .Y(N892) );
  AOI2BB2X1TF U1021 ( .B0(N2390), .B1(N695), .A0N(\GR[0][13] ), .A1N(N238), 
        .Y(N891) );
  AOI2BB2X1TF U1022 ( .B0(N2390), .B1(N696), .A0N(\GR[0][14] ), .A1N(N238), 
        .Y(N890) );
  AOI2BB2X1TF U1023 ( .B0(N2390), .B1(N697), .A0N(\GR[0][15] ), .A1N(N238), 
        .Y(N889) );
  AOI2BB2X1TF U1024 ( .B0(N233), .B1(N690), .A0N(N1363), .A1N(N232), .Y(N888)
         );
  AOI2BB2X1TF U1025 ( .B0(N233), .B1(N691), .A0N(N1362), .A1N(N232), .Y(N887)
         );
  AOI2BB2X1TF U1026 ( .B0(N233), .B1(N692), .A0N(N1361), .A1N(N232), .Y(N886)
         );
  AOI2BB2X1TF U1027 ( .B0(N233), .B1(N693), .A0N(N1360), .A1N(N232), .Y(N885)
         );
  AOI2BB2X1TF U1028 ( .B0(N233), .B1(N694), .A0N(N1359), .A1N(N232), .Y(N884)
         );
  AOI2BB2X1TF U1029 ( .B0(N233), .B1(N695), .A0N(N1358), .A1N(N232), .Y(N883)
         );
  AOI2BB2X1TF U1030 ( .B0(N233), .B1(N696), .A0N(N1357), .A1N(N232), .Y(N882)
         );
  AOI2BB2X1TF U1031 ( .B0(N233), .B1(N697), .A0N(N1356), .A1N(N232), .Y(N881)
         );
  AOI2BB2X1TF U1032 ( .B0(N229), .B1(N690), .A0N(N40), .A1N(N228), .Y(N880) );
  AOI2BB2X1TF U1033 ( .B0(N229), .B1(N691), .A0N(N41), .A1N(N229), .Y(N879) );
  AOI2BB2X1TF U1034 ( .B0(N229), .B1(N692), .A0N(N42), .A1N(N228), .Y(N878) );
  AOI2BB2X1TF U1035 ( .B0(N229), .B1(N693), .A0N(IO_DATAOUTA[11]), .A1N(N228), 
        .Y(N877) );
  AOI2BB2X1TF U1036 ( .B0(N229), .B1(N694), .A0N(N43), .A1N(N228), .Y(N876) );
  AOI2BB2X1TF U1037 ( .B0(N229), .B1(N695), .A0N(N1366), .A1N(N228), .Y(N875)
         );
  AOI2BB2X1TF U1038 ( .B0(N229), .B1(N696), .A0N(N1365), .A1N(N228), .Y(N874)
         );
  AOI2BB2X1TF U1039 ( .B0(N228), .B1(N697), .A0N(N1364), .A1N(N228), .Y(N873)
         );
  AOI2BB2X1TF U1040 ( .B0(N235), .B1(N690), .A0N(IO_DATAOUTB[8]), .A1N(N234), 
        .Y(N872) );
  AOI2BB2X1TF U1041 ( .B0(N235), .B1(N691), .A0N(IO_DATAOUTB[9]), .A1N(N234), 
        .Y(N871) );
  AOI2BB2X1TF U1042 ( .B0(N235), .B1(N692), .A0N(IO_DATAOUTB[10]), .A1N(N234), 
        .Y(N870) );
  AOI2BB2X1TF U1043 ( .B0(N235), .B1(N693), .A0N(N44), .A1N(N234), .Y(N869) );
  AOI2BB2X1TF U1044 ( .B0(N235), .B1(N694), .A0N(IO_DATAOUTB[12]), .A1N(N234), 
        .Y(N868) );
  AOI2BB2X1TF U1045 ( .B0(N235), .B1(N695), .A0N(N1369), .A1N(N234), .Y(N867)
         );
  AOI2BB2X1TF U1046 ( .B0(N235), .B1(N696), .A0N(N1368), .A1N(N234), .Y(N866)
         );
  AOI2BB2X1TF U1047 ( .B0(N235), .B1(N697), .A0N(N1367), .A1N(N234), .Y(N865)
         );
  AOI2BB2X1TF U1048 ( .B0(N237), .B1(N690), .A0N(IO_OFFSET[8]), .A1N(N236), 
        .Y(N864) );
  AOI2BB2X1TF U1049 ( .B0(N237), .B1(N691), .A0N(IO_OFFSET[9]), .A1N(N236), 
        .Y(N863) );
  AOI2BB2X1TF U1050 ( .B0(N237), .B1(N692), .A0N(N1375), .A1N(N236), .Y(N862)
         );
  AOI2BB2X1TF U1051 ( .B0(N237), .B1(N693), .A0N(N1374), .A1N(N236), .Y(N861)
         );
  AOI2BB2X1TF U1052 ( .B0(N237), .B1(N694), .A0N(N1373), .A1N(N236), .Y(N860)
         );
  AOI2BB2X1TF U1053 ( .B0(N237), .B1(N695), .A0N(N1372), .A1N(N236), .Y(N859)
         );
  AOI2BB2X1TF U1054 ( .B0(N237), .B1(N696), .A0N(N1371), .A1N(N236), .Y(N858)
         );
  AOI2BB2X1TF U1055 ( .B0(N237), .B1(N697), .A0N(N1370), .A1N(N236), .Y(N857)
         );
  AOI2BB2X1TF U1056 ( .B0(N295), .B1(N690), .A0N(\GR[5][8] ), .A1N(N685), .Y(
        N856) );
  AOI2BB2X1TF U1057 ( .B0(N295), .B1(N691), .A0N(\GR[5][9] ), .A1N(N685), .Y(
        N855) );
  AOI2BB2X1TF U1058 ( .B0(N295), .B1(N692), .A0N(\GR[5][10] ), .A1N(N685), .Y(
        N854) );
  AOI2BB2X1TF U1059 ( .B0(N295), .B1(N693), .A0N(\GR[5][11] ), .A1N(N685), .Y(
        N853) );
  AOI2BB2X1TF U1060 ( .B0(N295), .B1(N694), .A0N(\GR[5][12] ), .A1N(N685), .Y(
        N852) );
  AOI2BB2X1TF U1061 ( .B0(N295), .B1(N695), .A0N(\GR[5][13] ), .A1N(N685), .Y(
        N851) );
  AOI2BB2X1TF U1062 ( .B0(N295), .B1(N696), .A0N(\GR[5][14] ), .A1N(N685), .Y(
        N850) );
  AOI2BB2X1TF U1063 ( .B0(N295), .B1(N697), .A0N(\GR[5][15] ), .A1N(N685), .Y(
        N849) );
  AOI2BB2X1TF U1064 ( .B0(N294), .B1(N690), .A0N(\GR[6][8] ), .A1N(N687), .Y(
        N848) );
  AOI2BB2X1TF U1065 ( .B0(N294), .B1(N691), .A0N(\GR[6][9] ), .A1N(N687), .Y(
        N847) );
  AOI2BB2X1TF U1066 ( .B0(N294), .B1(N692), .A0N(\GR[6][10] ), .A1N(N687), .Y(
        N846) );
  AOI2BB2X1TF U1067 ( .B0(N294), .B1(N693), .A0N(\GR[6][11] ), .A1N(N687), .Y(
        N845) );
  AOI2BB2X1TF U1068 ( .B0(N294), .B1(N694), .A0N(\GR[6][12] ), .A1N(N687), .Y(
        N844) );
  AOI2BB2X1TF U1069 ( .B0(N294), .B1(N695), .A0N(\GR[6][13] ), .A1N(N687), .Y(
        N843) );
  AOI2BB2X1TF U1070 ( .B0(N294), .B1(N696), .A0N(\GR[6][14] ), .A1N(N687), .Y(
        N842) );
  AOI2BB2X1TF U1071 ( .B0(N294), .B1(N697), .A0N(\GR[6][15] ), .A1N(N687), .Y(
        N841) );
  AOI2BB2X1TF U1072 ( .B0(N231), .B1(N690), .A0N(\GR[7][8] ), .A1N(N230), .Y(
        N840) );
  AOI2BB2X1TF U1073 ( .B0(N231), .B1(N691), .A0N(\GR[7][9] ), .A1N(N230), .Y(
        N839) );
  AOI2BB2X1TF U1074 ( .B0(N231), .B1(N692), .A0N(\GR[7][10] ), .A1N(N230), .Y(
        N838) );
  AOI2BB2X1TF U1075 ( .B0(N231), .B1(N693), .A0N(\GR[7][11] ), .A1N(N230), .Y(
        N837) );
  AOI2BB2X1TF U1076 ( .B0(N231), .B1(N694), .A0N(\GR[7][12] ), .A1N(N230), .Y(
        N836) );
  AOI2BB2X1TF U1077 ( .B0(N231), .B1(N695), .A0N(\GR[7][13] ), .A1N(N230), .Y(
        N835) );
  AOI2BB2X1TF U1078 ( .B0(N231), .B1(N696), .A0N(\GR[7][14] ), .A1N(N230), .Y(
        N834) );
  AOI2BB2X1TF U1079 ( .B0(N231), .B1(N697), .A0N(\GR[7][15] ), .A1N(N230), .Y(
        N833) );
  NAND2X1TF U1080 ( .A(I_ADDR[2]), .B(I_ADDR[1]), .Y(N699) );
  XOR2X1TF U1081 ( .A(I_ADDR[5]), .B(N703), .Y(N704) );
  OAI2BB1X1TF U1082 ( .A0N(D_ADDR[5]), .A1N(N719), .B0(N705), .Y(N832) );
  NOR4XLTF U1083 ( .A(\IO_CONTROL[4] ), .B(\IO_CONTROL[5] ), .C(
        \IO_CONTROL[6] ), .D(\IO_CONTROL[7] ), .Y(N720) );
  NOR4XLTF U1084 ( .A(IO_STATUS[0]), .B(IO_STATUS[1]), .C(IO_STATUS[2]), .D(
        N720), .Y(N723) );
  NAND2X1TF U1085 ( .A(N734), .B(N1134), .Y(NEXT_STATE[2]) );
  NAND2X1TF U1087 ( .A(N302), .B(REG_A[4]), .Y(N739) );
  NAND2X1TF U1088 ( .A(N747), .B(REG_A[5]), .Y(N759) );
  NAND2X1TF U1089 ( .A(N808), .B(REG_A[7]), .Y(N752) );
  NAND4X1TF U1090 ( .A(N739), .B(N738), .C(N759), .D(N752), .Y(N822) );
  NAND2X1TF U1091 ( .A(N747), .B(REG_A[9]), .Y(N754) );
  NAND2X1TF U1092 ( .A(N808), .B(REG_A[11]), .Y(N1034) );
  NAND4BX1TF U1093 ( .AN(N741), .B(N754), .C(N740), .D(N1034), .Y(N987) );
  AOI222XLTF U1094 ( .A0(N822), .A1(N1043), .B0(N987), .B1(N1009), .C0(N742), 
        .C1(N767), .Y(N746) );
  NAND2X1TF U1095 ( .A(N1030), .B(REG_A[9]), .Y(N811) );
  NAND2X1TF U1096 ( .A(N808), .B(REG_A[4]), .Y(N774) );
  NAND2X1TF U1097 ( .A(N1031), .B(REG_A[7]), .Y(N812) );
  NAND2X1TF U1098 ( .A(REG_A[2]), .B(N747), .Y(N773) );
  OAI221XLTF U1099 ( .A0(N198), .A1(REG_A[14]), .B0(N354), .B1(REG_A[15]), 
        .C0(N355), .Y(N971) );
  NAND2X1TF U1100 ( .A(N1019), .B(N751), .Y(N795) );
  NAND2X1TF U1101 ( .A(N2130), .B(REG_A[8]), .Y(N788) );
  NAND4X1TF U1102 ( .A(N754), .B(N753), .C(N752), .D(N788), .Y(N1042) );
  NAND2X1TF U1103 ( .A(N613), .B(N1009), .Y(N983) );
  NAND2X1TF U1104 ( .A(N1031), .B(REG_A[6]), .Y(N789) );
  OAI222X1TF U1105 ( .A0(N829), .A1(N1016), .B0(N991), .B1(N1038), .C0(N995), 
        .C1(N1036), .Y(N772) );
  OAI221XLTF U1106 ( .A0(REG_A[1]), .A1(N357), .B0(N332), .B1(N1013), .C0(N376), .Y(N781) );
  NAND2X1TF U1107 ( .A(REG_A[3]), .B(N1030), .Y(N775) );
  NAND2X1TF U1108 ( .A(N778), .B(N356), .Y(N997) );
  NAND4BX1TF U1109 ( .AN(N791), .B(N790), .C(N789), .D(N788), .Y(N969) );
  NAND3X1TF U1110 ( .A(N804), .B(N803), .C(N802), .Y(N428) );
  NAND2X1TF U1111 ( .A(N1019), .B(N1009), .Y(N979) );
  NAND4BX1TF U1112 ( .AN(N814), .B(N813), .C(N812), .D(N811), .Y(N978) );
  AO21X1TF U1113 ( .A0(N360), .A1(N388), .B0(N815), .Y(N818) );
  NAND2X1TF U1114 ( .A(N1031), .B(REG_A[15]), .Y(N1015) );
  AOI2BB2X1TF U1115 ( .B0(REG_A[3]), .B1(N818), .A0N(N360), .A1N(N817), .Y(
        N819) );
  OAI2BB2XLTF U1116 ( .B0(N1039), .B1(N973), .A0N(N1009), .A1N(N1045), .Y(N974) );
  AOI2BB2X1TF U1117 ( .B0(N492), .B1(N268), .A0N(N992), .A1N(N991), .Y(N1002)
         );
  AOI222XLTF U1118 ( .A0(N1012), .A1(N1046), .B0(N1011), .B1(N1043), .C0(N1010), .C1(N1009), .Y(N1021) );
  AOI2BB2X1TF U1119 ( .B0(N239), .B1(N222), .A0N(N1085), .A1N(N572), .Y(N1070)
         );
  OAI31X1TF U1120 ( .A0(N1100), .A1(N1099), .A2(N1098), .B0(N1104), .Y(N1108)
         );
  AO22X1TF U1121 ( .A0(N1134), .A1(N372), .B0(N1133), .B1(I_DATAIN[7]), .Y(
        N507) );
  AO22X1TF U1122 ( .A0(N1134), .A1(N94), .B0(N1133), .B1(I_DATAIN[6]), .Y(N508) );
  AO22X1TF U1123 ( .A0(N1134), .A1(N93), .B0(N1133), .B1(I_DATAIN[5]), .Y(N509) );
  AO22X1TF U1124 ( .A0(N1134), .A1(N92), .B0(N1133), .B1(I_DATAIN[4]), .Y(N510) );
  AO22X1TF U1125 ( .A0(N1134), .A1(N97), .B0(N1133), .B1(I_DATAIN[2]), .Y(N512) );
  AO22X1TF U1126 ( .A0(N1134), .A1(N96), .B0(N1133), .B1(I_DATAIN[1]), .Y(N513) );
  AO22X1TF U1127 ( .A0(N1134), .A1(N95), .B0(N1133), .B1(I_DATAIN[0]), .Y(N514) );
  AO22X1TF U1128 ( .A0(N1139), .A1(N29), .B0(N1138), .B1(I_DATAIN[7]), .Y(N517) );
  AO22X1TF U1129 ( .A0(N1139), .A1(CODE_TYPE[3]), .B0(N1138), .B1(I_DATAIN[6]), 
        .Y(N518) );
  AO22X1TF U1130 ( .A0(N1139), .A1(N2000), .B0(N1138), .B1(I_DATAIN[5]), .Y(
        N519) );
  AO22X1TF U1131 ( .A0(N1139), .A1(N307), .B0(N1138), .B1(I_DATAIN[4]), .Y(
        N520) );
  AO22X1TF U1132 ( .A0(N1139), .A1(N91), .B0(N1138), .B1(I_DATAIN[2]), .Y(N522) );
  AO22X1TF U1133 ( .A0(N1139), .A1(N90), .B0(N1138), .B1(I_DATAIN[1]), .Y(N523) );
  AO22X1TF U1134 ( .A0(N1139), .A1(N89), .B0(N1138), .B1(I_DATAIN[0]), .Y(N524) );
  NAND4X1TF U1135 ( .A(N1148), .B(N1149), .C(N1150), .D(N1151), .Y(N177) );
  NAND4X1TF U1136 ( .A(N1152), .B(N1153), .C(N1154), .D(N1155), .Y(N176) );
  NAND4X1TF U1137 ( .A(N1156), .B(N1157), .C(N1158), .D(N1159), .Y(N175) );
  NAND4X1TF U1138 ( .A(N1160), .B(N1161), .C(N1162), .D(N1163), .Y(N174) );
  NAND4X1TF U1139 ( .A(N1164), .B(N1165), .C(N1166), .D(N1167), .Y(N173) );
  NAND4X1TF U1140 ( .A(N1168), .B(N1169), .C(N1170), .D(N1171), .Y(N172) );
  NAND4X1TF U1141 ( .A(N1172), .B(N1173), .C(N1174), .D(N1175), .Y(N171) );
  NAND4X1TF U1142 ( .A(N1176), .B(N1177), .C(N1178), .D(N1179), .Y(N170) );
  NAND4X1TF U1143 ( .A(N1180), .B(N1181), .C(N1182), .D(N1183), .Y(N169) );
  NAND4X1TF U1144 ( .A(N1184), .B(N1185), .C(N1186), .D(N1187), .Y(N168) );
  NAND4X1TF U1145 ( .A(N1188), .B(N1189), .C(N1190), .D(N1191), .Y(N167) );
  NAND4X1TF U1146 ( .A(N1192), .B(N1193), .C(N1194), .D(N1195), .Y(N166) );
  NAND4X1TF U1147 ( .A(N1196), .B(N1197), .C(N1198), .D(N1199), .Y(N165) );
  NAND4X1TF U1148 ( .A(N1200), .B(N1201), .C(N1202), .D(N1203), .Y(N164) );
  NAND4X1TF U1149 ( .A(N1204), .B(N1205), .C(N1206), .D(N1207), .Y(N163) );
  NAND4X1TF U1150 ( .A(N1208), .B(N1209), .C(N1210), .D(N1211), .Y(N162) );
  NAND4X1TF U1151 ( .A(N1220), .B(N1221), .C(N1222), .D(N1223), .Y(N214) );
  NAND4X1TF U1152 ( .A(N1224), .B(N1225), .C(N1226), .D(N1227), .Y(N213) );
  NAND4X1TF U1153 ( .A(N1228), .B(N1229), .C(N1230), .D(N1231), .Y(N212) );
  NAND4X1TF U1154 ( .A(N1232), .B(N1233), .C(N1234), .D(N1235), .Y(N211) );
  NAND4X1TF U1155 ( .A(N1236), .B(N1237), .C(N1238), .D(N1239), .Y(N210) );
  NAND4X1TF U1156 ( .A(N1240), .B(N1241), .C(N1242), .D(N1243), .Y(N209) );
  NAND4X1TF U1157 ( .A(N1244), .B(N1245), .C(N1246), .D(N1247), .Y(N208) );
  NAND4X1TF U1158 ( .A(N1248), .B(N1249), .C(N1250), .D(N1251), .Y(N207) );
  NAND4X1TF U1159 ( .A(N1252), .B(N1253), .C(N1254), .D(N1255), .Y(N206) );
  NAND4X1TF U1160 ( .A(N1256), .B(N1257), .C(N1258), .D(N1259), .Y(N205) );
  NAND4X1TF U1161 ( .A(N1260), .B(N1261), .C(N1262), .D(N1263), .Y(N204) );
  NAND4X1TF U1162 ( .A(N1264), .B(N1265), .C(N1266), .D(N1267), .Y(N203) );
  NAND4X1TF U1163 ( .A(N1268), .B(N1269), .C(N1270), .D(N1271), .Y(N202) );
  NAND4X1TF U1164 ( .A(N1272), .B(N1273), .C(N1274), .D(N1275), .Y(N201) );
  NAND4X1TF U1165 ( .A(N1276), .B(N1277), .C(N1278), .D(N1279), .Y(N200) );
  NAND4X1TF U1166 ( .A(N1280), .B(N1281), .C(N1282), .D(N1283), .Y(N199) );
  NAND4X1TF U1167 ( .A(N1292), .B(N1293), .C(N1294), .D(N1295), .Y(N254) );
  NAND4X1TF U1168 ( .A(N1296), .B(N1297), .C(N1298), .D(N1299), .Y(N253) );
  NAND4X1TF U1169 ( .A(N1300), .B(N1301), .C(N1302), .D(N1303), .Y(N252) );
  NAND4X1TF U1170 ( .A(N1304), .B(N1305), .C(N1306), .D(N1307), .Y(N251) );
  NAND4X1TF U1171 ( .A(N1308), .B(N1309), .C(N1310), .D(N1311), .Y(N250) );
  NAND4X1TF U1172 ( .A(N1312), .B(N1313), .C(N1314), .D(N1315), .Y(N249) );
  NAND4X1TF U1173 ( .A(N1316), .B(N1317), .C(N1318), .D(N1319), .Y(N248) );
  NAND4X1TF U1174 ( .A(N1320), .B(N1321), .C(N1322), .D(N1323), .Y(N247) );
  NAND4X1TF U1175 ( .A(N1324), .B(N1325), .C(N1326), .D(N1327), .Y(N246) );
  NAND4X1TF U1176 ( .A(N1328), .B(N1329), .C(N1330), .D(N1331), .Y(N245) );
  NAND4X1TF U1177 ( .A(N1332), .B(N1333), .C(N1334), .D(N1335), .Y(N244) );
  NAND4X1TF U1178 ( .A(N1336), .B(N1337), .C(N1338), .D(N1339), .Y(N243) );
  NAND4X1TF U1179 ( .A(N1340), .B(N1341), .C(N1342), .D(N1343), .Y(N242) );
  NAND4X1TF U1180 ( .A(N1344), .B(N1345), .C(N1346), .D(N1347), .Y(N241) );
  NAND4X1TF U1181 ( .A(N1348), .B(N1349), .C(N1350), .D(N1351), .Y(N240) );
  NAND4X1TF U1182 ( .A(N1352), .B(N1353), .C(N1354), .D(N1355), .Y(N239) );
endmodule


module SCPU_SRAM_8BIT_ALU_SPI_TOP_VG ( CLK, RST_N, CTRL_MODE, CTRL_BGN, CPU_BGN, 
        LOAD_N, CTRL_SI, APP_DONE, ADC_PI, TEST_MUX, CPU_WAIT, CTRL_RDY, 
        APP_START, CTRL_SO, NXT, SCLK1, SCLK2, LAT, SPI_SO );
  input [1:0] CTRL_MODE;
  input [9:0] ADC_PI;
  input [2:0] TEST_MUX;
  output [1:0] NXT;
  input CLK, RST_N, CTRL_BGN, CPU_BGN, LOAD_N, CTRL_SI, APP_DONE, CPU_WAIT;
  output CTRL_RDY, APP_START, CTRL_SO, SCLK1, SCLK2, LAT, SPI_SO;
  wire   CEN_AFTER_MUX, WEN_AFTER_MUX, I_CLK, I_RST_N, I_CTRL_BGN, I_CPU_BGN,
         I_LOAD_N, I_CTRL_SI, I_APP_DONE, I_CPU_WAIT, I_APP_START, I_CTRL_SO,
         I_SCLK1, I_SCLK2, I_LAT, I_SPI_SO, SCPU_CTRL_SPI_I_SPI_SO,
         \SCPU_CTRL_SPI_POUT[0] , \SCPU_CTRL_SPI_POUT[1] ,
         \SCPU_CTRL_SPI_POUT[2] , \SCPU_CTRL_SPI_POUT[3] ,
         \SCPU_CTRL_SPI_POUT[4] , \SCPU_CTRL_SPI_POUT[5] ,
         \SCPU_CTRL_SPI_POUT[6] , \SCPU_CTRL_SPI_POUT[7] ,
         \SCPU_CTRL_SPI_POUT[8] , \SCPU_CTRL_SPI_POUT[9] ,
         \SCPU_CTRL_SPI_POUT[10] , \SCPU_CTRL_SPI_POUT[11] ,
         \SCPU_CTRL_SPI_POUT[12] , \SCPU_CTRL_SPI_FOUT[0] ,
         \SCPU_CTRL_SPI_FOUT[1] , \SCPU_CTRL_SPI_FOUT[2] ,
         \SCPU_CTRL_SPI_FOUT[3] , \SCPU_CTRL_SPI_FOUT[4] ,
         \SCPU_CTRL_SPI_FOUT[5] , \SCPU_CTRL_SPI_FOUT[6] ,
         \SCPU_CTRL_SPI_FOUT[7] , \SCPU_CTRL_SPI_FOUT[8] ,
         \SCPU_CTRL_SPI_FOUT[9] , \SCPU_CTRL_SPI_FOUT[10] ,
         \SCPU_CTRL_SPI_FOUT[11] , \SCPU_CTRL_SPI_FOUT[12] , SCPU_CTRL_SPI_CEN,
         \SCPU_CTRL_SPI_IO_DATAOUTB[0] , \SCPU_CTRL_SPI_IO_DATAOUTB[1] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[2] , \SCPU_CTRL_SPI_IO_DATAOUTB[3] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[4] , \SCPU_CTRL_SPI_IO_DATAOUTB[5] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[6] , \SCPU_CTRL_SPI_IO_DATAOUTB[7] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[8] , \SCPU_CTRL_SPI_IO_DATAOUTB[9] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[10] , \SCPU_CTRL_SPI_IO_DATAOUTB[11] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[12] , \SCPU_CTRL_SPI_IO_DATAOUTA[0] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[1] , \SCPU_CTRL_SPI_IO_DATAOUTA[2] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[3] , \SCPU_CTRL_SPI_IO_DATAOUTA[4] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[5] , \SCPU_CTRL_SPI_IO_DATAOUTA[6] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[7] , \SCPU_CTRL_SPI_IO_DATAOUTA[8] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[9] , \SCPU_CTRL_SPI_IO_DATAOUTA[10] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[11] , \SCPU_CTRL_SPI_IO_DATAOUTA[12] ,
         \SCPU_CTRL_SPI_IO_DATAINA[0] , \SCPU_CTRL_SPI_IO_DATAINA[1] ,
         \SCPU_CTRL_SPI_IO_DATAINA[2] , \SCPU_CTRL_SPI_IO_DATAINA[3] ,
         \SCPU_CTRL_SPI_IO_DATAINA[4] , \SCPU_CTRL_SPI_IO_DATAINA[5] ,
         \SCPU_CTRL_SPI_IO_DATAINA[6] , \SCPU_CTRL_SPI_IO_DATAINA[7] ,
         \SCPU_CTRL_SPI_IO_DATAINA[8] , \SCPU_CTRL_SPI_IO_DATAINA[9] ,
         \SCPU_CTRL_SPI_IO_DATAINA[10] , \SCPU_CTRL_SPI_IO_DATAINA[11] ,
         \SCPU_CTRL_SPI_IO_DATAINA[12] , SCPU_CTRL_SPI_IO_CONTROL_0,
         SCPU_CTRL_SPI_IO_CONTROL_1, SCPU_CTRL_SPI_IO_CONTROL_2,
         SCPU_CTRL_SPI_IO_CONTROL_3, SCPU_CTRL_SPI_IO_CONTROL_4,
         SCPU_CTRL_SPI_IO_CONTROL_5, SCPU_CTRL_SPI_IO_CONTROL_6,
         \SCPU_CTRL_SPI_IO_STATUS[0] , SCPU_CTRL_SPI_D_WE,
         SCPU_CTRL_SPI_IS_I_ADDR, SCPU_CTRL_SPI_CCT_N57, SCPU_CTRL_SPI_CCT_N56,
         SCPU_CTRL_SPI_CCT_N55, SCPU_CTRL_SPI_CCT_N53, SCPU_CTRL_SPI_CCT_N52,
         SCPU_CTRL_SPI_CCT_IS_SHIFT, \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[3] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[5] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[7] , \SCPU_CTRL_SPI_CCT_REG_BITS[1] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[2] , \SCPU_CTRL_SPI_CCT_REG_BITS[3] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[4] , \SCPU_CTRL_SPI_CCT_REG_BITS[5] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[6] , \SCPU_CTRL_SPI_CCT_REG_BITS[7] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[8] , \SCPU_CTRL_SPI_CCT_REG_BITS[9] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[10] , \SCPU_CTRL_SPI_CCT_REG_BITS[11] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[12] , \SCPU_CTRL_SPI_CCT_REG_BITS[13] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[14] , \SCPU_CTRL_SPI_CCT_REG_BITS[15] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[16] , \SCPU_CTRL_SPI_CCT_REG_BITS[17] ,
         \SCPU_CTRL_SPI_CCT_CTRL_STATE[0] , SCPU_CTRL_SPI_PUT_N112,
         SCPU_CTRL_SPI_PUT_N111, SCPU_CTRL_SPI_PUT_N110,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] , SCPU_CTRL_SPI_PUT_N27,
         SCPU_CTRL_SPI_PUT_IS_ADDR_LEN_NZ, \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ,
         \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ,
         \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] ,
         \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[4] , \SCPU_CTRL_SPI_PUT_SPI_STATE[1] ,
         \SCPU_CTRL_SPI_PUT_CNT_STATE[0] , \SCPU_CTRL_SPI_PUT_CNT_STATE[1] ,
         \SCPU_CTRL_SPI_PUT_CNT_STATE[2] , N34, N35, N36, N37, N38, N39, N40,
         N41, N42, N43, N44, N45, N46, N47, N48, N87, N88, N89, N90, N91, N92,
         N93, N94, N95, N96, N100, N102, N108, N110, N111, N168, N174, N175,
         N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243,
         N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254,
         N256, N257, N258, N259, N260, N261, N263, N264, N265, N266, N277,
         N278, N279, N280, N281, N309, N310, N311, N312, N313, N314, N315,
         N316, N317, N318, N321, N322, N323, N324, N325, N326, N327, N328,
         N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, N339,
         N340, N341, N342, N343, N344, N345, N346, N347, N348, N349, N350,
         N351, N352, N353, N354, N355, N356, N357, N358, N359, N360, N361,
         N362, N363, N364, N365, N366, N367, N368, N369, N370, N371, N372,
         N373, N374, N375, N376, N377, N378, N379, N380, N381, N382, N383,
         N384, N385, N386, N387, N388, N389, N390, N391, N392, N393, N394,
         N395, N396, N397, N398, N399, N400, N401, N402, N403, N404, N405,
         N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416,
         N417, N418, N419, N420, N421, N422, N423, N424, N425, N426, N427,
         N428, N429, N430, N431, N432, N433, N434, N435, N436, N437, N438,
         N439, N440, N441, N442, N443, N444, N445, N446, N447, N448, N449,
         N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460,
         N461, N462, N463, N464, N465, N466, N467, N468, N469, N470, N471,
         N472, N473, N474, N475, N476, N477, N478, N479, N480, N481, N482,
         N483, N484, N485, N486, N487, N488, N489, N490, N491, N492, N493,
         N494, N495, N496, N497, N498, N499, N500, N501, N502, N503, N504,
         N505, N506, N507, N508, N509, N510, N511, N512, N513, N514, N515,
         N516;
  wire   [9:0] A_AFTER_MUX;
  wire   [7:0] D_AFTER_MUX;
  wire   [7:0] Q_FROM_SRAM;
  wire   [1:0] I_CTRL_MODE;
  wire   [9:0] I_ADC_PI;
  wire   [2:0] I_TEST_MUX;
  wire   [1:0] I_NXT;
  wire   [9:0] SCPU_CTRL_SPI_A_SPI;
  wire   [9:0] SCPU_CTRL_SPI_IO_OFFSET;
  wire   [7:0] SCPU_CTRL_SPI_D_DATAOUT;
  wire   [9:1] SCPU_CTRL_SPI_D_ADDR;
  wire   [9:0] SCPU_CTRL_SPI_I_ADDR;
  wire   [1:0] SCPU_CTRL_SPI_I_NXT;
  wire   [7:0] SCPU_CTRL_SPI_D_DATAIN;
  wire   [7:0] SCPU_CTRL_SPI_I_DATAIN;
  wire   [7:1] SCPU_CTRL_SPI_PUT_SRAM_REGS;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12;

  RA1SHD_IBM1024X8 sram ( .Q(Q_FROM_SRAM), .A(A_AFTER_MUX), .D(D_AFTER_MUX), 
        .CLK(I_CLK), .CEN(CEN_AFTER_MUX), .WEN(WEN_AFTER_MUX) );
  PIC ipad_clk ( .IE(1'b1), .P(CLK), .Y(I_CLK) );
  PIC ipad_rst_n ( .IE(1'b1), .P(RST_N), .Y(I_RST_N) );
  PIC ipad_ctrl_mode0 ( .IE(1'b1), .P(CTRL_MODE[0]), .Y(I_CTRL_MODE[0]) );
  PIC ipad_ctrl_mode1 ( .IE(1'b1), .P(CTRL_MODE[1]), .Y(I_CTRL_MODE[1]) );
  PIC ipad_ctrl_bgn ( .IE(1'b1), .P(CTRL_BGN), .Y(I_CTRL_BGN) );
  PIC ipad_cpu_bgn ( .IE(1'b1), .P(CPU_BGN), .Y(I_CPU_BGN) );
  PIC ipad_load_n ( .IE(1'b1), .P(LOAD_N), .Y(I_LOAD_N) );
  PIC ipad_ctrl_si ( .IE(1'b1), .P(CTRL_SI), .Y(I_CTRL_SI) );
  PIC ipad_app_done ( .IE(1'b1), .P(APP_DONE), .Y(I_APP_DONE) );
  PIC ipad_adc_pi0 ( .IE(1'b1), .P(ADC_PI[0]), .Y(I_ADC_PI[0]) );
  PIC ipad_adc_pi1 ( .IE(1'b1), .P(ADC_PI[1]), .Y(I_ADC_PI[1]) );
  PIC ipad_adc_pi2 ( .IE(1'b1), .P(ADC_PI[2]), .Y(I_ADC_PI[2]) );
  PIC ipad_adc_pi3 ( .IE(1'b1), .P(ADC_PI[3]), .Y(I_ADC_PI[3]) );
  PIC ipad_adc_pi4 ( .IE(1'b1), .P(ADC_PI[4]), .Y(I_ADC_PI[4]) );
  PIC ipad_adc_pi5 ( .IE(1'b1), .P(ADC_PI[5]), .Y(I_ADC_PI[5]) );
  PIC ipad_adc_pi6 ( .IE(1'b1), .P(ADC_PI[6]), .Y(I_ADC_PI[6]) );
  PIC ipad_adc_pi7 ( .IE(1'b1), .P(ADC_PI[7]), .Y(I_ADC_PI[7]) );
  PIC ipad_adc_pi8 ( .IE(1'b1), .P(ADC_PI[8]), .Y(I_ADC_PI[8]) );
  PIC ipad_adc_pi9 ( .IE(1'b1), .P(ADC_PI[9]), .Y(I_ADC_PI[9]) );
  PIC ipad_test_mux0 ( .IE(1'b1), .P(TEST_MUX[0]), .Y(I_TEST_MUX[0]) );
  PIC ipad_test_mux1 ( .IE(1'b1), .P(TEST_MUX[1]), .Y(I_TEST_MUX[1]) );
  PIC ipad_test_mux2 ( .IE(1'b1), .P(TEST_MUX[2]), .Y(I_TEST_MUX[2]) );
  PIC ipad_cpu_wait ( .IE(1'b1), .P(CPU_WAIT), .Y(I_CPU_WAIT) );
  POC8B opad_app_start ( .A(I_APP_START), .P(APP_START) );
  POC8B opad_ctrl_rdy ( .A(N265), .P(CTRL_RDY) );
  POC8B opad_ctrl_so ( .A(I_CTRL_SO), .P(CTRL_SO) );
  POC8B opad_nxt0 ( .A(I_NXT[0]), .P(NXT[0]) );
  POC8B opad_nxt1 ( .A(I_NXT[1]), .P(NXT[1]) );
  POC8B opad_sclk1 ( .A(I_SCLK1), .P(SCLK1) );
  POC8B opad_sclk2 ( .A(I_SCLK2), .P(SCLK2) );
  POC8B opad_lat ( .A(I_LAT), .P(LAT) );
  POC8B opad_spi_so ( .A(I_SPI_SO), .P(SPI_SO) );
  SHARE_SUPERALU_VG \scpu_ctrl_spi/ALU_01  ( .CLK(I_CLK), .RST_N(I_RST_N), .X_IN(
        {\SCPU_CTRL_SPI_IO_DATAOUTA[12] , \SCPU_CTRL_SPI_IO_DATAOUTA[11] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[10] , \SCPU_CTRL_SPI_IO_DATAOUTA[9] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[8] , \SCPU_CTRL_SPI_IO_DATAOUTA[7] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[6] , \SCPU_CTRL_SPI_IO_DATAOUTA[5] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[4] , \SCPU_CTRL_SPI_IO_DATAOUTA[3] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[2] , \SCPU_CTRL_SPI_IO_DATAOUTA[1] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[0] }), .Y_IN({
        \SCPU_CTRL_SPI_IO_DATAOUTB[12] , \SCPU_CTRL_SPI_IO_DATAOUTB[11] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[10] , \SCPU_CTRL_SPI_IO_DATAOUTB[9] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[8] , \SCPU_CTRL_SPI_IO_DATAOUTB[7] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[6] , \SCPU_CTRL_SPI_IO_DATAOUTB[5] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[4] , \SCPU_CTRL_SPI_IO_DATAOUTB[3] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[2] , \SCPU_CTRL_SPI_IO_DATAOUTB[1] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[0] }), .ALU_START(N316), .ALU_TYPE({
        SCPU_CTRL_SPI_IO_CONTROL_4, SCPU_CTRL_SPI_IO_CONTROL_3, 
        SCPU_CTRL_SPI_IO_CONTROL_2}), .MODE_TYPE({SCPU_CTRL_SPI_IO_CONTROL_1, 
        SCPU_CTRL_SPI_IO_CONTROL_0}), .OFFSET(SCPU_CTRL_SPI_IO_OFFSET), .FOUT(
        {\SCPU_CTRL_SPI_FOUT[12] , \SCPU_CTRL_SPI_FOUT[11] , 
        \SCPU_CTRL_SPI_FOUT[10] , \SCPU_CTRL_SPI_FOUT[9] , 
        \SCPU_CTRL_SPI_FOUT[8] , \SCPU_CTRL_SPI_FOUT[7] , 
        \SCPU_CTRL_SPI_FOUT[6] , \SCPU_CTRL_SPI_FOUT[5] , 
        \SCPU_CTRL_SPI_FOUT[4] , \SCPU_CTRL_SPI_FOUT[3] , 
        \SCPU_CTRL_SPI_FOUT[2] , \SCPU_CTRL_SPI_FOUT[1] , 
        \SCPU_CTRL_SPI_FOUT[0] }), .POUT({\SCPU_CTRL_SPI_POUT[12] , 
        \SCPU_CTRL_SPI_POUT[11] , \SCPU_CTRL_SPI_POUT[10] , 
        \SCPU_CTRL_SPI_POUT[9] , \SCPU_CTRL_SPI_POUT[8] , 
        \SCPU_CTRL_SPI_POUT[7] , \SCPU_CTRL_SPI_POUT[6] , 
        \SCPU_CTRL_SPI_POUT[5] , \SCPU_CTRL_SPI_POUT[4] , 
        \SCPU_CTRL_SPI_POUT[3] , \SCPU_CTRL_SPI_POUT[2] , 
        \SCPU_CTRL_SPI_POUT[1] , \SCPU_CTRL_SPI_POUT[0] }), .ALU_IS_DONE(
        \SCPU_CTRL_SPI_IO_STATUS[0] ) );
  SERIAL_CPU_8BIT_VG \scpu_ctrl_spi/uut  ( .CLK(I_CLK), .ENABLE(1'b0), .RST_N(
        I_RST_N), .START(I_CPU_BGN), .I_DATAIN(SCPU_CTRL_SPI_I_DATAIN), 
        .D_DATAIN(SCPU_CTRL_SPI_D_DATAIN), .CPU_WAIT(I_CPU_WAIT), .IS_I_ADDR(
        SCPU_CTRL_SPI_IS_I_ADDR), .NXT(SCPU_CTRL_SPI_I_NXT), .I_ADDR(
        SCPU_CTRL_SPI_I_ADDR), .D_ADDR({SCPU_CTRL_SPI_D_ADDR, 
        SYNOPSYS_UNCONNECTED__0}), .D_WE(SCPU_CTRL_SPI_D_WE), .D_DATAOUT(
        SCPU_CTRL_SPI_D_DATAOUT), .IO_STATUS({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, I_APP_DONE, N266, 
        \SCPU_CTRL_SPI_IO_STATUS[0] }), .IO_DATAINA({1'b0, 1'b0, 1'b0, 
        \SCPU_CTRL_SPI_IO_DATAINA[12] , \SCPU_CTRL_SPI_IO_DATAINA[11] , 
        \SCPU_CTRL_SPI_IO_DATAINA[10] , \SCPU_CTRL_SPI_IO_DATAINA[9] , 
        \SCPU_CTRL_SPI_IO_DATAINA[8] , \SCPU_CTRL_SPI_IO_DATAINA[7] , 
        \SCPU_CTRL_SPI_IO_DATAINA[6] , \SCPU_CTRL_SPI_IO_DATAINA[5] , 
        \SCPU_CTRL_SPI_IO_DATAINA[4] , \SCPU_CTRL_SPI_IO_DATAINA[3] , 
        \SCPU_CTRL_SPI_IO_DATAINA[2] , \SCPU_CTRL_SPI_IO_DATAINA[1] , 
        \SCPU_CTRL_SPI_IO_DATAINA[0] }), .IO_DATAINB({1'b0, 1'b0, 1'b0, 
        \SCPU_CTRL_SPI_POUT[12] , \SCPU_CTRL_SPI_POUT[11] , 
        \SCPU_CTRL_SPI_POUT[10] , \SCPU_CTRL_SPI_POUT[9] , 
        \SCPU_CTRL_SPI_POUT[8] , \SCPU_CTRL_SPI_POUT[7] , 
        \SCPU_CTRL_SPI_POUT[6] , \SCPU_CTRL_SPI_POUT[5] , 
        \SCPU_CTRL_SPI_POUT[4] , \SCPU_CTRL_SPI_POUT[3] , 
        \SCPU_CTRL_SPI_POUT[2] , \SCPU_CTRL_SPI_POUT[1] , 
        \SCPU_CTRL_SPI_POUT[0] }), .IO_DATAOUTA({SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        \SCPU_CTRL_SPI_IO_DATAOUTA[12] , \SCPU_CTRL_SPI_IO_DATAOUTA[11] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[10] , \SCPU_CTRL_SPI_IO_DATAOUTA[9] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[8] , \SCPU_CTRL_SPI_IO_DATAOUTA[7] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[6] , \SCPU_CTRL_SPI_IO_DATAOUTA[5] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[4] , \SCPU_CTRL_SPI_IO_DATAOUTA[3] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[2] , \SCPU_CTRL_SPI_IO_DATAOUTA[1] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[0] }), .IO_DATAOUTB({
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, \SCPU_CTRL_SPI_IO_DATAOUTB[12] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[11] , \SCPU_CTRL_SPI_IO_DATAOUTB[10] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[9] , \SCPU_CTRL_SPI_IO_DATAOUTB[8] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[7] , \SCPU_CTRL_SPI_IO_DATAOUTB[6] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[5] , \SCPU_CTRL_SPI_IO_DATAOUTB[4] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[3] , \SCPU_CTRL_SPI_IO_DATAOUTB[2] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[1] , \SCPU_CTRL_SPI_IO_DATAOUTB[0] }), 
        .IO_OFFSET({SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SCPU_CTRL_SPI_IO_OFFSET}), .\IO_CONTROL[7] (I_APP_START), 
        .\IO_CONTROL[6] (SCPU_CTRL_SPI_IO_CONTROL_6), .\IO_CONTROL[5]_BAR (
        SCPU_CTRL_SPI_IO_CONTROL_5), .\IO_CONTROL[4] (
        SCPU_CTRL_SPI_IO_CONTROL_4), .\IO_CONTROL[3] (
        SCPU_CTRL_SPI_IO_CONTROL_3), .\IO_CONTROL[2] (
        SCPU_CTRL_SPI_IO_CONTROL_2), .\IO_CONTROL[1] (
        SCPU_CTRL_SPI_IO_CONTROL_1), .\IO_CONTROL[0] (
        SCPU_CTRL_SPI_IO_CONTROL_0) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[7]  ( .D(N168), .RN(
        SCPU_CTRL_SPI_CCT_N57), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[7] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[5]  ( .D(N168), .RN(
        SCPU_CTRL_SPI_CCT_N55), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[5] ), .QN(N333) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[3]  ( .D(N168), .RN(
        SCPU_CTRL_SPI_CCT_N53), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[3] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[2]  ( .D(N168), .RN(
        SCPU_CTRL_SPI_CCT_N52), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ), .QN(N335) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[6]  ( .D(N168), .RN(
        SCPU_CTRL_SPI_CCT_N56), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[17]  ( .D(I_CTRL_SI), .E(N342), 
        .CK(I_CLK), .Q(\SCPU_CTRL_SPI_CCT_REG_BITS[17] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[16]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[17] ), .E(N342), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[16] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[15]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[16] ), .E(N100), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[15] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[14]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[15] ), .E(N100), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[14] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[13]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[14] ), .E(N100), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[13] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[12]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[13] ), .E(N100), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[12] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[11]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[12] ), .E(N100), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[11] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[10]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[11] ), .E(N100), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[10] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[9]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[10] ), .E(N100), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[9] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[8]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[9] ), .E(N100), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[8] ) );
  DFFSX2TF \scpu_ctrl_spi/put/cnt_state_reg[0]  ( .D(SCPU_CTRL_SPI_PUT_N110), 
        .CK(I_CLK), .SN(SCPU_CTRL_SPI_IO_CONTROL_6), .Q(
        \SCPU_CTRL_SPI_PUT_CNT_STATE[0] ), .QN(N334) );
  DFFRX2TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[3]  ( .D(N252), .CK(I_CLK), 
        .RN(N315), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ), .QN(N338) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[2]  ( .D(N42), .CK(I_CLK), 
        .SN(N41), .RN(N40), .QN(N337) );
  DFFRX2TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[0]  ( .D(N249), .CK(I_CLK), 
        .RN(N315), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .QN(N332) );
  DFFRX2TF \scpu_ctrl_spi/put/spi_state_reg[0]  ( .D(N253), .CK(I_CLK), .RN(
        N315), .Q(N328), .QN(N108) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[4]  ( .D(N48), .CK(I_CLK), 
        .SN(N47), .RN(N46), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[4] ), .QN(N326)
         );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[1]  ( .D(N39), .CK(I_CLK), 
        .SN(N38), .RN(N37), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ), .QN(N324)
         );
  DFFRX2TF \scpu_ctrl_spi/put/cnt_state_reg[1]  ( .D(SCPU_CTRL_SPI_PUT_N111), 
        .CK(I_CLK), .RN(N315), .Q(\SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .QN(N323)
         );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[3]  ( .D(N45), .CK(I_CLK), 
        .SN(N44), .RN(N43), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] ), .QN(N322)
         );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[7]  ( .D(N248), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[7]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[6]  ( .D(N242), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[6]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[5]  ( .D(N243), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[5]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[4]  ( .D(N244), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[4]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[3]  ( .D(N245), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[3]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[2]  ( .D(N246), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[2]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[1]  ( .D(N247), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[1]) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[7]  ( .D(N233), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[7] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[6]  ( .D(N234), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[6] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[5]  ( .D(N235), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[5] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[4]  ( .D(N236), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[4] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[3]  ( .D(N237), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[3] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[2]  ( .D(N238), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[2] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[1]  ( .D(N239), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[1] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/is_shift_reg  ( .D(N174), .RN(N175), .CK(I_CLK), 
        .QN(SCPU_CTRL_SPI_CCT_IS_SHIFT) );
  DFFQX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[1]  ( .D(N258), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[4]  ( .D(N260), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[0]  ( .D(N259), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[0]  ( .D(N240), .CK(I_CLK), .Q(
        I_CTRL_SO) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[0]  ( .D(N241), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_I_SPI_SO) );
  DFFXLTF \scpu_ctrl_spi/cct/ctrl_state_reg[0]  ( .D(N261), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .QN(N339) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[0]  ( .D(N36), .CK(I_CLK), 
        .SN(N35), .RN(N34), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ) );
  DFFRX2TF \scpu_ctrl_spi/put/spi_state_reg[2]  ( .D(N256), .CK(I_CLK), .RN(
        N315), .Q(N321), .QN(N110) );
  DFFNSRX4TF \scpu_ctrl_spi/put/spi_MUX_reg  ( .D(N257), .CKN(I_CLK), .SN(1'b1), .RN(1'b1), .Q(N340), .QN(N111) );
  DFFNSRXLTF \scpu_ctrl_spi/cct/CEN_reg  ( .D(N264), .CKN(I_CLK), .SN(1'b1), 
        .RN(1'b1), .Q(SCPU_CTRL_SPI_CEN) );
  DFFNSRXLTF \scpu_ctrl_spi/put/is_addr_len_nz_reg  ( .D(SCPU_CTRL_SPI_PUT_N27), .CKN(I_CLK), .SN(1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_PUT_IS_ADDR_LEN_NZ) );
  DFFNSRXLTF \scpu_ctrl_spi/put/sram_addr_reg[9]  ( .D(N96), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[9]) );
  EDFFTRXLTF \scpu_ctrl_spi/cct/ctrl_state_reg[1]  ( .RN(I_CTRL_BGN), .D(1'b1), 
        .E(N281), .CK(I_CLK), .Q(N325), .QN(N102) );
  DFFRX1TF \scpu_ctrl_spi/put/cnt_state_reg[2]  ( .D(SCPU_CTRL_SPI_PUT_N112), 
        .CK(I_CLK), .RN(N315), .Q(\SCPU_CTRL_SPI_PUT_CNT_STATE[2] ) );
  DFFRX1TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[1]  ( .D(N250), .CK(I_CLK), 
        .RN(N315), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ) );
  DFFRX1TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[2]  ( .D(N251), .CK(I_CLK), 
        .RN(N314), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ) );
  DFFRX2TF \scpu_ctrl_spi/put/spi_state_reg[1]  ( .D(N254), .CK(I_CLK), .RN(
        N315), .Q(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[1]  ( .D(N88), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[1]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[3]  ( .D(N90), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[3]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[2]  ( .D(N89), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[2]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[6]  ( .D(N93), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[6]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[4]  ( .D(N91), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[4]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[7]  ( .D(N94), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[7]), .QN(N329) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[8]  ( .D(N95), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[8]), .QN(N331) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[0]  ( .D(N87), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[0]), .QN(N330) );
  DFFNSRX2TF \scpu_ctrl_spi/cct/D_WE_reg  ( .D(N263), .CKN(I_CLK), .SN(1'b1), 
        .RN(1'b1), .QN(N327) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[5]  ( .D(N92), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[5]), .QN(N336) );
  NOR3BX2TF U290 ( .AN(N337), .B(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .C(
        \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ), .Y(N515) );
  INVX2TF U291 ( .A(SCPU_CTRL_SPI_IO_CONTROL_5), .Y(N309) );
  AND2X2TF U292 ( .A(N311), .B(N327), .Y(N370) );
  AOI22XLTF U293 ( .A0(SCPU_CTRL_SPI_A_SPI[8]), .A1(N365), .B0(
        SCPU_CTRL_SPI_I_ADDR[8]), .B1(N364), .Y(N277) );
  AOI22XLTF U294 ( .A0(SCPU_CTRL_SPI_D_ADDR[8]), .A1(N366), .B0(N310), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[16] ), .Y(N278) );
  NAND2X1TF U295 ( .A(N277), .B(N278), .Y(A_AFTER_MUX[8]) );
  OAI22X1TF U296 ( .A0(SCPU_CTRL_SPI_PUT_IS_ADDR_LEN_NZ), .A1(N511), .B0(N423), 
        .B1(N321), .Y(N279) );
  AOI21X1TF U297 ( .A0(N423), .A1(N321), .B0(N279), .Y(N280) );
  AOI22X1TF U298 ( .A0(N425), .A1(N280), .B0(N110), .B1(N428), .Y(N256) );
  OA21XLTF U299 ( .A0(N317), .A1(I_CTRL_MODE[0]), .B0(N410), .Y(N281) );
  AOI22XLTF U300 ( .A0(SCPU_CTRL_SPI_A_SPI[3]), .A1(N365), .B0(
        SCPU_CTRL_SPI_I_ADDR[3]), .B1(N364), .Y(N355) );
  AOI22XLTF U301 ( .A0(SCPU_CTRL_SPI_A_SPI[1]), .A1(N365), .B0(
        SCPU_CTRL_SPI_I_ADDR[1]), .B1(N364), .Y(N351) );
  AOI22XLTF U302 ( .A0(N366), .A1(SCPU_CTRL_SPI_D_ADDR[9]), .B0(N310), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[17] ), .Y(N367) );
  OR2X2TF U318 ( .A(SCPU_CTRL_SPI_CEN), .B(N439), .Y(N369) );
  INVX2TF U319 ( .A(I_TEST_MUX[1]), .Y(N374) );
  NAND2XLTF U320 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[3] ), .B(N345), .Y(N44) );
  NAND2XLTF U321 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[4] ), .B(N345), .Y(N47) );
  NAND2BXLTF U322 ( .AN(\SCPU_CTRL_SPI_IO_DATAOUTB[2] ), .B(N341), .Y(N40) );
  NAND2XLTF U323 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[1] ), .B(N345), .Y(N38) );
  NAND2XLTF U324 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[2] ), .B(N345), .Y(N41) );
  NAND2BXLTF U325 ( .AN(\SCPU_CTRL_SPI_IO_DATAOUTB[1] ), .B(N341), .Y(N37) );
  NAND2XLTF U326 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[0] ), .B(N345), .Y(N35) );
  NAND2BXLTF U327 ( .AN(\SCPU_CTRL_SPI_IO_DATAOUTB[0] ), .B(N345), .Y(N34) );
  NAND2BXLTF U328 ( .AN(\SCPU_CTRL_SPI_IO_DATAOUTB[3] ), .B(N341), .Y(N43) );
  NAND2BXLTF U329 ( .AN(\SCPU_CTRL_SPI_IO_DATAOUTB[4] ), .B(N341), .Y(N46) );
  AOI22X1TF U330 ( .A0(SCPU_CTRL_SPI_D_ADDR[3]), .A1(N366), .B0(N310), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[11] ), .Y(N354) );
  OAI211XLTF U331 ( .A0(N427), .A1(N328), .B0(N321), .C0(N425), .Y(N426) );
  AND3X2TF U332 ( .A(N314), .B(N516), .C(SCPU_CTRL_SPI_PUT_IS_ADDR_LEN_NZ), 
        .Y(N507) );
  INVX2TF U333 ( .A(N341), .Y(N314) );
  NAND2XLTF U334 ( .A(SCPU_CTRL_SPI_A_SPI[0]), .B(SCPU_CTRL_SPI_A_SPI[1]), .Y(
        N504) );
  INVX2TF U335 ( .A(SCPU_CTRL_SPI_IO_CONTROL_6), .Y(N341) );
  CLKBUFX2TF U336 ( .A(\SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .Y(N317) );
  INVX2TF U337 ( .A(N369), .Y(N310) );
  INVX2TF U338 ( .A(N369), .Y(N311) );
  INVX2TF U339 ( .A(N507), .Y(N312) );
  INVX2TF U340 ( .A(N507), .Y(N313) );
  INVX2TF U341 ( .A(N341), .Y(N315) );
  INVX2TF U342 ( .A(SCPU_CTRL_SPI_IO_CONTROL_5), .Y(N316) );
  OAI211X1TF U343 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] ), .A1(
        \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[4] ), .B0(N516), .C0(N515), .Y(N514)
         );
  NAND4BX2TF U344 ( .AN(N264), .B(I_CTRL_BGN), .C(SCPU_CTRL_SPI_CCT_IS_SHIFT), 
        .D(N453), .Y(N463) );
  AOI32XLTF U345 ( .A0(N516), .A1(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] ), .A2(
        N515), .B0(N514), .B1(N322), .Y(N45) );
  NOR3X4TF U346 ( .A(N108), .B(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .C(N321), 
        .Y(N516) );
  INVX2TF U347 ( .A(I_CTRL_BGN), .Y(N318) );
  NOR3X4TF U348 ( .A(N441), .B(N440), .C(N344), .Y(N450) );
  AOI32X1TF U349 ( .A0(N111), .A1(N439), .A2(SCPU_CTRL_SPI_D_WE), .B0(
        I_CTRL_BGN), .B1(N327), .Y(WEN_AFTER_MUX) );
  INVX2TF U350 ( .A(I_CTRL_BGN), .Y(N439) );
  NAND4X1TF U351 ( .A(N397), .B(N396), .C(N395), .D(N394), .Y(I_SCLK2) );
  NOR2X1TF U352 ( .A(N427), .B(N442), .Y(N438) );
  NOR3XLTF U353 ( .A(N317), .B(N325), .C(N439), .Y(N414) );
  NAND2X1TF U354 ( .A(I_CTRL_BGN), .B(N413), .Y(N420) );
  NOR2X1TF U355 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[3] ), .B(N346), .Y(N174)
         );
  CLKBUFX2TF U356 ( .A(N100), .Y(N342) );
  NAND2X1TF U357 ( .A(N361), .B(N360), .Y(A_AFTER_MUX[6]) );
  NAND2X1TF U358 ( .A(N359), .B(N358), .Y(A_AFTER_MUX[5]) );
  NAND2X1TF U359 ( .A(N357), .B(N356), .Y(A_AFTER_MUX[4]) );
  NAND2X1TF U360 ( .A(N355), .B(N354), .Y(A_AFTER_MUX[3]) );
  NAND2X1TF U361 ( .A(N353), .B(N352), .Y(A_AFTER_MUX[2]) );
  NAND2X1TF U362 ( .A(N351), .B(N350), .Y(A_AFTER_MUX[1]) );
  NAND2X1TF U363 ( .A(N368), .B(N367), .Y(A_AFTER_MUX[9]) );
  NAND2X1TF U364 ( .A(N363), .B(N362), .Y(A_AFTER_MUX[7]) );
  NOR2X2TF U365 ( .A(N340), .B(N464), .Y(N366) );
  NOR2X2TF U366 ( .A(N340), .B(N472), .Y(N364) );
  CLKBUFX2TF U367 ( .A(N509), .Y(N343) );
  NAND4X1TF U368 ( .A(N379), .B(N378), .C(N377), .D(N376), .Y(I_LAT) );
  NAND4X1TF U369 ( .A(N387), .B(N386), .C(N385), .D(N384), .Y(I_NXT[1]) );
  NAND4X1TF U370 ( .A(N383), .B(N382), .C(N381), .D(N380), .Y(I_NXT[0]) );
  NAND4X1TF U371 ( .A(N409), .B(N408), .C(N407), .D(N406), .Y(I_SPI_SO) );
  NAND4X1TF U372 ( .A(N392), .B(N391), .C(N390), .D(N389), .Y(I_SCLK1) );
  AO22X1TF U373 ( .A0(N316), .A1(\SCPU_CTRL_SPI_FOUT[4] ), .B0(N474), .B1(
        I_ADC_PI[4]), .Y(\SCPU_CTRL_SPI_IO_DATAINA[4] ) );
  AO22X1TF U374 ( .A0(N309), .A1(\SCPU_CTRL_SPI_FOUT[3] ), .B0(N474), .B1(
        I_ADC_PI[3]), .Y(\SCPU_CTRL_SPI_IO_DATAINA[3] ) );
  INVX2TF U375 ( .A(I_TEST_MUX[0]), .Y(N373) );
  INVX2TF U376 ( .A(I_TEST_MUX[2]), .Y(N372) );
  AO21X1TF U377 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[3] ), .A1(N346), .B0(
        N174), .Y(SCPU_CTRL_SPI_CCT_N53) );
  OAI2BB2XLTF U378 ( .B0(N478), .B1(N477), .A0N(
        \SCPU_CTRL_SPI_PUT_CNT_STATE[2] ), .A1N(N476), .Y(
        SCPU_CTRL_SPI_PUT_N112) );
  NAND2X1TF U379 ( .A(N516), .B(N510), .Y(N512) );
  NOR2X1TF U380 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ), .B(N347), .Y(N348)
         );
  NAND2X1TF U381 ( .A(N333), .B(N411), .Y(N347) );
  NOR2X1TF U382 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ), .B(N412), .Y(N411)
         );
  NAND2X1TF U383 ( .A(N174), .B(N175), .Y(N413) );
  OR3X1TF U384 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ), .B(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .C(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ), .Y(N346) );
  NAND3X1TF U385 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .B(N110), .C(N328), 
        .Y(N437) );
  AND3X2TF U386 ( .A(SCPU_CTRL_SPI_CCT_IS_SHIFT), .B(N102), .C(N317), .Y(N100)
         );
  OAI2BB2XLTF U387 ( .B0(N428), .B1(N479), .A0N(
        \SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .A1N(N426), .Y(N254) );
  NOR2X1TF U388 ( .A(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ), .B(N424), .Y(N427)
         );
  OAI2BB1X1TF U389 ( .A0N(N311), .A1N(\SCPU_CTRL_SPI_CCT_REG_BITS[8] ), .B0(
        N349), .Y(A_AFTER_MUX[0]) );
  AO22X1TF U390 ( .A0(N370), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[7] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[7]), .B1(N439), .Y(D_AFTER_MUX[7]) );
  AO22X1TF U391 ( .A0(N370), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[6] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[6]), .B1(N439), .Y(D_AFTER_MUX[6]) );
  AO22X1TF U392 ( .A0(N370), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[5] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[5]), .B1(N439), .Y(D_AFTER_MUX[5]) );
  AO22X1TF U393 ( .A0(N370), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[4] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[4]), .B1(N318), .Y(D_AFTER_MUX[4]) );
  AO22X1TF U394 ( .A0(N370), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[3] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[3]), .B1(N318), .Y(D_AFTER_MUX[3]) );
  AO22X1TF U395 ( .A0(N370), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[2] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[2]), .B1(N318), .Y(D_AFTER_MUX[2]) );
  AO22X1TF U396 ( .A0(N370), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[1] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[1]), .B1(N318), .Y(D_AFTER_MUX[1]) );
  AO22X1TF U397 ( .A0(N370), .A1(I_CTRL_SO), .B0(SCPU_CTRL_SPI_D_DATAOUT[0]), 
        .B1(N318), .Y(D_AFTER_MUX[0]) );
  NAND2X2TF U398 ( .A(SCPU_CTRL_SPI_IS_I_ADDR), .B(N439), .Y(N472) );
  NOR2X2TF U399 ( .A(I_CTRL_BGN), .B(N111), .Y(N365) );
  NAND2X1TF U400 ( .A(N317), .B(N325), .Y(N264) );
  NAND2BX2TF U401 ( .AN(SCPU_CTRL_SPI_IS_I_ADDR), .B(N439), .Y(N464) );
  CLKBUFX2TF U402 ( .A(N341), .Y(N345) );
  CLKBUFX2TF U403 ( .A(N341), .Y(N344) );
  NAND2X1TF U404 ( .A(N516), .B(SCPU_CTRL_SPI_PUT_IS_ADDR_LEN_NZ), .Y(N479) );
  INVX2TF U405 ( .A(N309), .Y(N474) );
  OAI21X1TF U406 ( .A0(N418), .A1(N335), .B0(N346), .Y(SCPU_CTRL_SPI_CCT_N52)
         );
  NOR2X1TF U407 ( .A(\SCPU_CTRL_SPI_PUT_CNT_STATE[0] ), .B(N475), .Y(
        SCPU_CTRL_SPI_PUT_N110) );
  OAI211X1TF U408 ( .A0(N438), .A1(N332), .B0(N437), .C0(N436), .Y(N249) );
  AOI31X1TF U409 ( .A0(N516), .A1(N515), .A2(N322), .B0(N326), .Y(N48) );
  OAI211X1TF U410 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .A1(N436), .B0(
        N437), .C0(N435), .Y(N250) );
  OAI21X1TF U411 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .A1(N478), .B0(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .Y(N435) );
  OAI31X1TF U412 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .A1(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .A2(N478), .B0(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ), .Y(N434) );
  AOI22X1TF U413 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ), .A1(N432), .B0(
        N433), .B1(N338), .Y(N252) );
  AOI21X1TF U414 ( .A0(N440), .A1(N424), .B0(N478), .Y(N432) );
  NOR2X1TF U415 ( .A(N441), .B(N438), .Y(N478) );
  OAI21X1TF U416 ( .A0(N411), .A1(N333), .B0(N347), .Y(SCPU_CTRL_SPI_CCT_N55)
         );
  OAI32X1TF U417 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ), .A1(
        \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .A2(N512), .B0(N513), .B1(N324), 
        .Y(N39) );
  AOI32X1TF U418 ( .A0(N513), .A1(N514), .A2(N324), .B0(N337), .B1(N514), .Y(
        N42) );
  NOR2X1TF U419 ( .A(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .B(N511), .Y(N513)
         );
  OAI22X1TF U420 ( .A0(I_CTRL_MODE[1]), .A1(N417), .B0(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .B1(N420), .Y(N259) );
  OAI21X1TF U421 ( .A0(N415), .A1(N420), .B0(N419), .Y(N260) );
  AOI21X1TF U422 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ), .A1(N412), .B0(
        N411), .Y(N415) );
  INVX2TF U423 ( .A(N174), .Y(N412) );
  OAI21X1TF U424 ( .A0(N421), .A1(N420), .B0(N419), .Y(N258) );
  NOR3BX1TF U425 ( .AN(N414), .B(I_LOAD_N), .C(N413), .Y(N416) );
  AOI21X1TF U426 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .A1(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ), .B0(N418), .Y(N421) );
  NOR2X1TF U427 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ), .B(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .Y(N418) );
  INVX2TF U428 ( .A(N420), .Y(N168) );
  NOR4X1TF U429 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[7] ), .B(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ), .C(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[5] ), .D(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ), .Y(N175) );
  OAI21X1TF U430 ( .A0(N452), .A1(N471), .B0(N448), .Y(N242) );
  AOI22X1TF U431 ( .A0(N450), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[6]), .B0(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[7]), .B1(N449), .Y(N448) );
  OAI21X1TF U432 ( .A0(N470), .A1(N452), .B0(N447), .Y(N243) );
  AOI22X1TF U433 ( .A0(N450), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[5]), .B0(N449), 
        .B1(SCPU_CTRL_SPI_PUT_SRAM_REGS[6]), .Y(N447) );
  OAI21X1TF U434 ( .A0(N469), .A1(N452), .B0(N446), .Y(N244) );
  AOI22X1TF U435 ( .A0(N450), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[4]), .B0(N449), 
        .B1(SCPU_CTRL_SPI_PUT_SRAM_REGS[5]), .Y(N446) );
  OAI21X1TF U436 ( .A0(N467), .A1(N452), .B0(N444), .Y(N246) );
  AOI22X1TF U437 ( .A0(N450), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[2]), .B0(N449), 
        .B1(SCPU_CTRL_SPI_PUT_SRAM_REGS[3]), .Y(N444) );
  OAI21X1TF U438 ( .A0(N465), .A1(N452), .B0(N451), .Y(N241) );
  AOI22X1TF U439 ( .A0(SCPU_CTRL_SPI_I_SPI_SO), .A1(N450), .B0(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[1]), .B1(N449), .Y(N451) );
  OAI21X1TF U440 ( .A0(N468), .A1(N452), .B0(N445), .Y(N245) );
  AOI22X1TF U441 ( .A0(N450), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[3]), .B0(N449), 
        .B1(SCPU_CTRL_SPI_PUT_SRAM_REGS[4]), .Y(N445) );
  OAI21X1TF U442 ( .A0(N466), .A1(N452), .B0(N443), .Y(N247) );
  AOI22X1TF U443 ( .A0(N450), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[1]), .B0(N449), 
        .B1(SCPU_CTRL_SPI_PUT_SRAM_REGS[2]), .Y(N443) );
  NOR2X2TF U444 ( .A(N344), .B(N442), .Y(N449) );
  INVX2TF U445 ( .A(N442), .Y(N440) );
  NAND3X2TF U446 ( .A(N439), .B(N315), .C(N441), .Y(N452) );
  INVX2TF U447 ( .A(N437), .Y(N441) );
  OAI21X1TF U448 ( .A0(N465), .A1(N463), .B0(N454), .Y(N240) );
  AOI22X1TF U449 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[1] ), .A1(N342), .B0(
        I_CTRL_SO), .B1(N461), .Y(N454) );
  OAI21X1TF U450 ( .A0(N468), .A1(N463), .B0(N457), .Y(N237) );
  AOI22X1TF U451 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[4] ), .A1(N342), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[3] ), .B1(N461), .Y(N457) );
  OAI21X1TF U452 ( .A0(N466), .A1(N463), .B0(N455), .Y(N239) );
  AOI22X1TF U453 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[2] ), .A1(N342), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[1] ), .B1(N461), .Y(N455) );
  OAI21X1TF U454 ( .A0(N473), .A1(N463), .B0(N462), .Y(N233) );
  AOI22X1TF U455 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[8] ), .A1(N342), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[7] ), .B1(N461), .Y(N462) );
  OAI21X1TF U456 ( .A0(N469), .A1(N463), .B0(N458), .Y(N236) );
  AOI22X1TF U457 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[5] ), .A1(N342), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[4] ), .B1(N461), .Y(N458) );
  OAI21X1TF U458 ( .A0(N467), .A1(N463), .B0(N456), .Y(N238) );
  AOI22X1TF U459 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[3] ), .A1(N342), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[2] ), .B1(N461), .Y(N456) );
  OAI21X1TF U460 ( .A0(N471), .A1(N463), .B0(N460), .Y(N234) );
  AOI22X1TF U461 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[7] ), .A1(N342), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[6] ), .B1(N461), .Y(N460) );
  OAI21X1TF U462 ( .A0(N470), .A1(N463), .B0(N459), .Y(N235) );
  AOI22X1TF U463 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[6] ), .A1(N342), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[5] ), .B1(N461), .Y(N459) );
  OAI211X4TF U464 ( .A0(N102), .A1(N453), .B0(N317), .C0(
        SCPU_CTRL_SPI_CCT_IS_SHIFT), .Y(N461) );
  INVX2TF U465 ( .A(I_CTRL_MODE[1]), .Y(N453) );
  NOR2X1TF U466 ( .A(N102), .B(N317), .Y(N265) );
  AND2X2TF U467 ( .A(SCPU_CTRL_SPI_CEN), .B(I_CTRL_BGN), .Y(CEN_AFTER_MUX) );
  AOI32X1TF U468 ( .A0(N430), .A1(N429), .A2(N479), .B0(N428), .B1(N429), .Y(
        N253) );
  OAI21X1TF U469 ( .A0(N321), .A1(N477), .B0(N328), .Y(N429) );
  INVX2TF U470 ( .A(N475), .Y(N477) );
  INVX2TF U471 ( .A(N428), .Y(N425) );
  INVX2TF U472 ( .A(N431), .Y(N424) );
  NOR3X1TF U473 ( .A(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ), .B(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .C(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .Y(N431) );
  AOI21X1TF U474 ( .A0(N321), .A1(N423), .B0(N475), .Y(N428) );
  NOR3X1TF U475 ( .A(\SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .B(
        \SCPU_CTRL_SPI_PUT_CNT_STATE[0] ), .C(\SCPU_CTRL_SPI_PUT_CNT_STATE[2] ), .Y(N475) );
  NOR2X1TF U476 ( .A(N473), .B(N472), .Y(SCPU_CTRL_SPI_I_DATAIN[7]) );
  NOR2X1TF U477 ( .A(N470), .B(N472), .Y(SCPU_CTRL_SPI_I_DATAIN[5]) );
  NOR2X1TF U478 ( .A(N466), .B(N472), .Y(SCPU_CTRL_SPI_I_DATAIN[1]) );
  NOR2X1TF U479 ( .A(N467), .B(N472), .Y(SCPU_CTRL_SPI_I_DATAIN[2]) );
  NOR2X1TF U480 ( .A(N471), .B(N472), .Y(SCPU_CTRL_SPI_I_DATAIN[6]) );
  NOR2X1TF U481 ( .A(N465), .B(N472), .Y(SCPU_CTRL_SPI_I_DATAIN[0]) );
  NOR2X1TF U482 ( .A(N469), .B(N472), .Y(SCPU_CTRL_SPI_I_DATAIN[4]) );
  NOR2X1TF U483 ( .A(N468), .B(N472), .Y(SCPU_CTRL_SPI_I_DATAIN[3]) );
  AND2X2TF U484 ( .A(N510), .B(N315), .Y(SCPU_CTRL_SPI_PUT_N27) );
  AOI22X1TF U485 ( .A0(SCPU_CTRL_SPI_D_ADDR[6]), .A1(N366), .B0(N310), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[14] ), .Y(N360) );
  AOI22X1TF U486 ( .A0(SCPU_CTRL_SPI_A_SPI[6]), .A1(N365), .B0(
        SCPU_CTRL_SPI_I_ADDR[6]), .B1(N364), .Y(N361) );
  AOI22X1TF U487 ( .A0(SCPU_CTRL_SPI_D_ADDR[5]), .A1(N366), .B0(N311), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[13] ), .Y(N358) );
  AOI22X1TF U488 ( .A0(SCPU_CTRL_SPI_A_SPI[5]), .A1(N365), .B0(
        SCPU_CTRL_SPI_I_ADDR[5]), .B1(N364), .Y(N359) );
  AOI22X1TF U489 ( .A0(SCPU_CTRL_SPI_D_ADDR[4]), .A1(N366), .B0(N311), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[12] ), .Y(N356) );
  AOI22X1TF U490 ( .A0(SCPU_CTRL_SPI_A_SPI[4]), .A1(N365), .B0(
        SCPU_CTRL_SPI_I_ADDR[4]), .B1(N364), .Y(N357) );
  AOI22X1TF U491 ( .A0(SCPU_CTRL_SPI_D_ADDR[2]), .A1(N366), .B0(N311), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[10] ), .Y(N352) );
  AOI22X1TF U492 ( .A0(SCPU_CTRL_SPI_A_SPI[2]), .A1(N365), .B0(
        SCPU_CTRL_SPI_I_ADDR[2]), .B1(N364), .Y(N353) );
  AOI22X1TF U493 ( .A0(SCPU_CTRL_SPI_D_ADDR[1]), .A1(N366), .B0(N311), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[9] ), .Y(N350) );
  AOI22X1TF U494 ( .A0(SCPU_CTRL_SPI_A_SPI[9]), .A1(N365), .B0(N364), .B1(
        SCPU_CTRL_SPI_I_ADDR[9]), .Y(N368) );
  AOI22X1TF U495 ( .A0(N366), .A1(SCPU_CTRL_SPI_D_ADDR[7]), .B0(N310), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[15] ), .Y(N362) );
  AOI22X1TF U496 ( .A0(SCPU_CTRL_SPI_A_SPI[7]), .A1(N365), .B0(N364), .B1(
        SCPU_CTRL_SPI_I_ADDR[7]), .Y(N363) );
  NOR2X1TF U497 ( .A(N467), .B(N464), .Y(SCPU_CTRL_SPI_D_DATAIN[2]) );
  NOR2X1TF U498 ( .A(N469), .B(N464), .Y(SCPU_CTRL_SPI_D_DATAIN[4]) );
  NOR2X1TF U499 ( .A(N471), .B(N464), .Y(SCPU_CTRL_SPI_D_DATAIN[6]) );
  NOR2X1TF U500 ( .A(N468), .B(N464), .Y(SCPU_CTRL_SPI_D_DATAIN[3]) );
  NOR2X1TF U501 ( .A(N465), .B(N464), .Y(SCPU_CTRL_SPI_D_DATAIN[0]) );
  NOR2X1TF U502 ( .A(N466), .B(N464), .Y(SCPU_CTRL_SPI_D_DATAIN[1]) );
  NOR2X1TF U503 ( .A(N473), .B(N464), .Y(SCPU_CTRL_SPI_D_DATAIN[7]) );
  NOR2X1TF U504 ( .A(N470), .B(N464), .Y(SCPU_CTRL_SPI_D_DATAIN[5]) );
  OAI32X1TF U505 ( .A0(N344), .A1(N111), .A2(N422), .B0(N511), .B1(N344), .Y(
        N257) );
  INVX2TF U506 ( .A(N516), .Y(N511) );
  NOR2X1TF U507 ( .A(N108), .B(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .Y(N422) );
  OAI21X1TF U508 ( .A0(N343), .A1(N330), .B0(N508), .Y(N87) );
  AOI22X1TF U509 ( .A0(N507), .A1(N330), .B0(\SCPU_CTRL_SPI_IO_DATAOUTA[0] ), 
        .B1(N344), .Y(N508) );
  AOI22X1TF U510 ( .A0(N486), .A1(N329), .B0(\SCPU_CTRL_SPI_IO_DATAOUTA[7] ), 
        .B1(N345), .Y(N487) );
  OAI21X1TF U511 ( .A0(SCPU_CTRL_SPI_A_SPI[5]), .A1(N494), .B0(N493), .Y(N92)
         );
  AOI22X1TF U512 ( .A0(SCPU_CTRL_SPI_A_SPI[5]), .A1(N492), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[5] ), .B1(N345), .Y(N493) );
  OAI21X1TF U513 ( .A0(N491), .A1(N313), .B0(N343), .Y(N492) );
  OAI31X1TF U514 ( .A0(SCPU_CTRL_SPI_A_SPI[3]), .A1(N313), .A2(N501), .B0(N500), .Y(N90) );
  AOI22X1TF U515 ( .A0(SCPU_CTRL_SPI_A_SPI[3]), .A1(N499), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[3] ), .B1(N344), .Y(N500) );
  OAI21X1TF U516 ( .A0(N498), .A1(N312), .B0(N343), .Y(N499) );
  OAI31X1TF U517 ( .A0(SCPU_CTRL_SPI_A_SPI[1]), .A1(N313), .A2(N330), .B0(N506), .Y(N88) );
  AOI22X1TF U518 ( .A0(SCPU_CTRL_SPI_A_SPI[1]), .A1(N505), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[1] ), .B1(N344), .Y(N506) );
  OAI21X1TF U519 ( .A0(SCPU_CTRL_SPI_A_SPI[0]), .A1(N312), .B0(N343), .Y(N505)
         );
  OAI31X1TF U520 ( .A0(SCPU_CTRL_SPI_A_SPI[2]), .A1(N313), .A2(N504), .B0(N503), .Y(N89) );
  AOI22X1TF U521 ( .A0(SCPU_CTRL_SPI_A_SPI[2]), .A1(N502), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[2] ), .B1(N344), .Y(N503) );
  AOI32X1TF U522 ( .A0(SCPU_CTRL_SPI_A_SPI[0]), .A1(N343), .A2(
        SCPU_CTRL_SPI_A_SPI[1]), .B0(N313), .B1(N343), .Y(N502) );
  OAI31X1TF U523 ( .A0(SCPU_CTRL_SPI_A_SPI[4]), .A1(N313), .A2(N497), .B0(N496), .Y(N91) );
  AOI22X1TF U524 ( .A0(SCPU_CTRL_SPI_A_SPI[4]), .A1(N495), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[4] ), .B1(N345), .Y(N496) );
  AOI32X1TF U525 ( .A0(N498), .A1(N343), .A2(SCPU_CTRL_SPI_A_SPI[3]), .B0(N313), .B1(N343), .Y(N495) );
  OAI31X1TF U526 ( .A0(SCPU_CTRL_SPI_A_SPI[6]), .A1(N336), .A2(N494), .B0(N490), .Y(N93) );
  AOI22X1TF U527 ( .A0(SCPU_CTRL_SPI_A_SPI[6]), .A1(N489), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[6] ), .B1(N345), .Y(N490) );
  AOI32X1TF U528 ( .A0(N491), .A1(N343), .A2(SCPU_CTRL_SPI_A_SPI[5]), .B0(N313), .B1(N343), .Y(N489) );
  OAI21X1TF U529 ( .A0(N485), .A1(N331), .B0(N484), .Y(N95) );
  OAI31X1TF U530 ( .A0(SCPU_CTRL_SPI_A_SPI[9]), .A1(N331), .A2(N483), .B0(N482), .Y(N96) );
  AOI22X1TF U531 ( .A0(SCPU_CTRL_SPI_A_SPI[9]), .A1(N481), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[9] ), .B1(N344), .Y(N482) );
  OAI21X1TF U532 ( .A0(SCPU_CTRL_SPI_A_SPI[8]), .A1(N313), .B0(N485), .Y(N481)
         );
  AOI21X1TF U533 ( .A0(N507), .A1(N329), .B0(N488), .Y(N485) );
  NOR2X1TF U534 ( .A(N312), .B(N480), .Y(N486) );
  INVX2TF U535 ( .A(N501), .Y(N498) );
  AND2X2TF U536 ( .A(\SCPU_CTRL_SPI_FOUT[11] ), .B(N309), .Y(
        \SCPU_CTRL_SPI_IO_DATAINA[11] ) );
  AND2X2TF U537 ( .A(\SCPU_CTRL_SPI_FOUT[12] ), .B(N309), .Y(
        \SCPU_CTRL_SPI_IO_DATAINA[12] ) );
  AOI21X1TF U538 ( .A0(SCPU_CTRL_SPI_D_ADDR[2]), .A1(N404), .B0(N375), .Y(N376) );
  AOI22X1TF U539 ( .A0(N403), .A1(Q_FROM_SRAM[1]), .B0(N402), .B1(
        SCPU_CTRL_SPI_I_ADDR[2]), .Y(N377) );
  AOI22X1TF U540 ( .A0(N401), .A1(\SCPU_CTRL_SPI_IO_DATAINA[1] ), .B0(N400), 
        .B1(\SCPU_CTRL_SPI_POUT[1] ), .Y(N378) );
  AOI22X1TF U541 ( .A0(N399), .A1(N266), .B0(N398), .B1(
        \SCPU_CTRL_SPI_FOUT[1] ), .Y(N379) );
  AOI22X1TF U542 ( .A0(N402), .A1(SCPU_CTRL_SPI_I_ADDR[6]), .B0(N405), .B1(
        SCPU_CTRL_SPI_I_NXT[1]), .Y(N385) );
  AOI22X1TF U543 ( .A0(N400), .A1(\SCPU_CTRL_SPI_POUT[5] ), .B0(N403), .B1(
        Q_FROM_SRAM[5]), .Y(N386) );
  AOI22X1TF U544 ( .A0(N398), .A1(\SCPU_CTRL_SPI_FOUT[5] ), .B0(N401), .B1(
        \SCPU_CTRL_SPI_IO_DATAINA[5] ), .Y(N387) );
  AOI22X1TF U545 ( .A0(N402), .A1(SCPU_CTRL_SPI_I_ADDR[5]), .B0(N405), .B1(
        SCPU_CTRL_SPI_I_NXT[0]), .Y(N381) );
  AOI22X1TF U546 ( .A0(N400), .A1(\SCPU_CTRL_SPI_POUT[4] ), .B0(N403), .B1(
        Q_FROM_SRAM[4]), .Y(N382) );
  AOI22X1TF U547 ( .A0(N398), .A1(\SCPU_CTRL_SPI_FOUT[4] ), .B0(N401), .B1(
        \SCPU_CTRL_SPI_IO_DATAINA[4] ), .Y(N383) );
  AND2X2TF U548 ( .A(\SCPU_CTRL_SPI_FOUT[10] ), .B(N309), .Y(
        \SCPU_CTRL_SPI_IO_DATAINA[10] ) );
  NOR3X1TF U549 ( .A(N108), .B(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .C(N110), 
        .Y(N266) );
  AOI22X1TF U550 ( .A0(N405), .A1(SCPU_CTRL_SPI_I_SPI_SO), .B0(N404), .B1(
        SCPU_CTRL_SPI_D_ADDR[1]), .Y(N406) );
  AOI22X1TF U551 ( .A0(N403), .A1(Q_FROM_SRAM[0]), .B0(N402), .B1(
        SCPU_CTRL_SPI_I_ADDR[1]), .Y(N407) );
  AOI22X1TF U552 ( .A0(N401), .A1(\SCPU_CTRL_SPI_IO_DATAINA[0] ), .B0(N400), 
        .B1(\SCPU_CTRL_SPI_POUT[0] ), .Y(N408) );
  AOI22X1TF U553 ( .A0(N399), .A1(\SCPU_CTRL_SPI_IO_STATUS[0] ), .B0(N398), 
        .B1(\SCPU_CTRL_SPI_FOUT[0] ), .Y(N409) );
  AOI22X1TF U554 ( .A0(N403), .A1(Q_FROM_SRAM[3]), .B0(N402), .B1(
        SCPU_CTRL_SPI_I_ADDR[4]), .Y(N390) );
  AOI22X1TF U555 ( .A0(N400), .A1(\SCPU_CTRL_SPI_POUT[3] ), .B0(N404), .B1(
        SCPU_CTRL_SPI_D_ADDR[4]), .Y(N391) );
  AOI22X1TF U556 ( .A0(N398), .A1(\SCPU_CTRL_SPI_FOUT[3] ), .B0(N401), .B1(
        \SCPU_CTRL_SPI_IO_DATAINA[3] ), .Y(N392) );
  AOI22X1TF U557 ( .A0(SCPU_CTRL_SPI_D_ADDR[3]), .A1(N404), .B0(N393), .B1(
        N323), .Y(N394) );
  AND3X2TF U558 ( .A(N340), .B(\SCPU_CTRL_SPI_PUT_CNT_STATE[0] ), .C(N405), 
        .Y(N393) );
  INVX2TF U559 ( .A(N388), .Y(N405) );
  NOR3X2TF U560 ( .A(N374), .B(N373), .C(N372), .Y(N404) );
  AOI22X1TF U561 ( .A0(Q_FROM_SRAM[2]), .A1(N403), .B0(N402), .B1(
        SCPU_CTRL_SPI_I_ADDR[3]), .Y(N395) );
  NOR3X2TF U562 ( .A(I_TEST_MUX[0]), .B(N374), .C(N372), .Y(N402) );
  NOR2X2TF U563 ( .A(I_TEST_MUX[1]), .B(N371), .Y(N403) );
  AOI22X1TF U564 ( .A0(N401), .A1(\SCPU_CTRL_SPI_IO_DATAINA[2] ), .B0(N400), 
        .B1(\SCPU_CTRL_SPI_POUT[2] ), .Y(N396) );
  NOR3X2TF U565 ( .A(I_TEST_MUX[2]), .B(N373), .C(N374), .Y(N400) );
  NOR3X2TF U566 ( .A(I_TEST_MUX[0]), .B(I_TEST_MUX[2]), .C(N374), .Y(N401) );
  AOI22X1TF U567 ( .A0(N399), .A1(I_APP_DONE), .B0(N398), .B1(
        \SCPU_CTRL_SPI_FOUT[2] ), .Y(N397) );
  NOR3X2TF U568 ( .A(I_TEST_MUX[1]), .B(I_TEST_MUX[2]), .C(N373), .Y(N398) );
  NOR3X1TF U569 ( .A(I_TEST_MUX[1]), .B(I_TEST_MUX[0]), .C(N372), .Y(N399) );
  INVX2TF U570 ( .A(Q_FROM_SRAM[2]), .Y(N467) );
  INVX2TF U571 ( .A(Q_FROM_SRAM[4]), .Y(N469) );
  INVX2TF U572 ( .A(Q_FROM_SRAM[6]), .Y(N471) );
  INVX2TF U573 ( .A(Q_FROM_SRAM[3]), .Y(N468) );
  INVX2TF U574 ( .A(Q_FROM_SRAM[0]), .Y(N465) );
  INVX2TF U575 ( .A(Q_FROM_SRAM[1]), .Y(N466) );
  INVX2TF U576 ( .A(Q_FROM_SRAM[7]), .Y(N473) );
  INVX2TF U577 ( .A(Q_FROM_SRAM[5]), .Y(N470) );
  NAND2X1TF U578 ( .A(N314), .B(N479), .Y(N509) );
  AO21X1TF U579 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ), .A1(N347), .B0(
        N348), .Y(SCPU_CTRL_SPI_CCT_N56) );
  XOR2X1TF U580 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[7] ), .B(N348), .Y(
        SCPU_CTRL_SPI_CCT_N57) );
  OAI221XLTF U581 ( .A0(N111), .A1(SCPU_CTRL_SPI_A_SPI[0]), .B0(N340), .B1(
        SCPU_CTRL_SPI_I_ADDR[0]), .C0(N439), .Y(N349) );
  AO22X1TF U582 ( .A0(N309), .A1(\SCPU_CTRL_SPI_FOUT[1] ), .B0(N474), .B1(
        I_ADC_PI[1]), .Y(\SCPU_CTRL_SPI_IO_DATAINA[1] ) );
  NAND2X1TF U583 ( .A(I_TEST_MUX[0]), .B(I_TEST_MUX[2]), .Y(N371) );
  NAND3X1TF U584 ( .A(N374), .B(N373), .C(N372), .Y(N388) );
  NOR4XLTF U585 ( .A(N110), .B(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .C(N328), 
        .D(N388), .Y(N375) );
  NAND2X1TF U586 ( .A(N404), .B(SCPU_CTRL_SPI_D_ADDR[5]), .Y(N380) );
  AO22X1TF U587 ( .A0(N309), .A1(\SCPU_CTRL_SPI_FOUT[5] ), .B0(N474), .B1(
        I_ADC_PI[5]), .Y(\SCPU_CTRL_SPI_IO_DATAINA[5] ) );
  NAND2X1TF U588 ( .A(N404), .B(SCPU_CTRL_SPI_D_ADDR[6]), .Y(N384) );
  NAND2X1TF U589 ( .A(\SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .B(N393), .Y(N389) );
  AO22X1TF U590 ( .A0(N316), .A1(\SCPU_CTRL_SPI_FOUT[2] ), .B0(N474), .B1(
        I_ADC_PI[2]), .Y(\SCPU_CTRL_SPI_IO_DATAINA[2] ) );
  AO22X1TF U591 ( .A0(N309), .A1(\SCPU_CTRL_SPI_FOUT[0] ), .B0(N474), .B1(
        I_ADC_PI[0]), .Y(\SCPU_CTRL_SPI_IO_DATAINA[0] ) );
  NAND2BX1TF U592 ( .AN(N264), .B(I_CTRL_MODE[1]), .Y(N263) );
  OAI221XLTF U593 ( .A0(N317), .A1(I_LOAD_N), .B0(N339), .B1(N413), .C0(
        I_CTRL_BGN), .Y(N410) );
  AO22X1TF U594 ( .A0(N317), .A1(N168), .B0(N414), .B1(N410), .Y(N261) );
  NAND2BX1TF U595 ( .AN(I_CTRL_MODE[0]), .B(N416), .Y(N419) );
  NAND2X1TF U596 ( .A(I_CTRL_MODE[0]), .B(N416), .Y(N417) );
  NAND2X1TF U597 ( .A(N108), .B(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .Y(N423) );
  NAND3X1TF U598 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .B(N108), .C(N321), 
        .Y(N442) );
  AOI2BB2X1TF U599 ( .B0(N427), .B1(N321), .A0N(N328), .A1N(
        \SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .Y(N430) );
  NAND2X1TF U600 ( .A(N431), .B(N438), .Y(N433) );
  NAND3X1TF U601 ( .A(N437), .B(N434), .C(N433), .Y(N251) );
  NAND2X1TF U602 ( .A(N438), .B(N332), .Y(N436) );
  OAI2BB2XLTF U603 ( .B0(N473), .B1(N452), .A0N(N450), .A1N(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[7]), .Y(N248) );
  AO22X1TF U604 ( .A0(N309), .A1(\SCPU_CTRL_SPI_FOUT[6] ), .B0(N474), .B1(
        I_ADC_PI[6]), .Y(\SCPU_CTRL_SPI_IO_DATAINA[6] ) );
  AO22X1TF U605 ( .A0(N316), .A1(\SCPU_CTRL_SPI_FOUT[7] ), .B0(N474), .B1(
        I_ADC_PI[7]), .Y(\SCPU_CTRL_SPI_IO_DATAINA[7] ) );
  AO22X1TF U606 ( .A0(N316), .A1(\SCPU_CTRL_SPI_FOUT[8] ), .B0(N474), .B1(
        I_ADC_PI[8]), .Y(\SCPU_CTRL_SPI_IO_DATAINA[8] ) );
  AO22X1TF U607 ( .A0(N309), .A1(\SCPU_CTRL_SPI_FOUT[9] ), .B0(N474), .B1(
        I_ADC_PI[9]), .Y(\SCPU_CTRL_SPI_IO_DATAINA[9] ) );
  AO22X1TF U608 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .A1(
        \SCPU_CTRL_SPI_PUT_CNT_STATE[0] ), .B0(N323), .B1(
        SCPU_CTRL_SPI_PUT_N110), .Y(SCPU_CTRL_SPI_PUT_N111) );
  NAND2X1TF U609 ( .A(N323), .B(N334), .Y(N476) );
  NAND3X1TF U610 ( .A(N326), .B(N322), .C(N515), .Y(N510) );
  NAND3X1TF U611 ( .A(SCPU_CTRL_SPI_A_SPI[2]), .B(SCPU_CTRL_SPI_A_SPI[0]), .C(
        SCPU_CTRL_SPI_A_SPI[1]), .Y(N501) );
  NAND2X1TF U612 ( .A(N498), .B(SCPU_CTRL_SPI_A_SPI[3]), .Y(N497) );
  NOR2BX1TF U613 ( .AN(SCPU_CTRL_SPI_A_SPI[4]), .B(N497), .Y(N491) );
  NAND3X1TF U614 ( .A(N491), .B(SCPU_CTRL_SPI_A_SPI[5]), .C(
        SCPU_CTRL_SPI_A_SPI[6]), .Y(N480) );
  NAND2X1TF U615 ( .A(SCPU_CTRL_SPI_A_SPI[7]), .B(N486), .Y(N483) );
  OAI2BB1X1TF U616 ( .A0N(N480), .A1N(N507), .B0(N509), .Y(N488) );
  AOI2BB2X1TF U617 ( .B0(\SCPU_CTRL_SPI_IO_DATAOUTA[8] ), .B1(N344), .A0N(
        SCPU_CTRL_SPI_A_SPI[8]), .A1N(N483), .Y(N484) );
  OAI2BB1X1TF U618 ( .A0N(SCPU_CTRL_SPI_A_SPI[7]), .A1N(N488), .B0(N487), .Y(
        N94) );
  NAND2X1TF U619 ( .A(N507), .B(N491), .Y(N494) );
  XNOR2X1TF U621 ( .A(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .B(N512), .Y(N36)
         );
endmodule

