
module SHARE_SUPERALU_VG ( CLK, RST_N, X_IN, Y_IN, ALU_START, ALU_TYPE, MODE_TYPE, 
        OFFSET, FOUT, POUT, ALU_IS_DONE );
  input [12:0] X_IN;
  input [12:0] Y_IN;
  input [2:0] ALU_TYPE;
  input [1:0] MODE_TYPE;
  input [9:0] OFFSET;
  output [12:0] FOUT;
  output [12:0] POUT;
  input CLK, RST_N, ALU_START;
  output ALU_IS_DONE;
  wire   POST_WORK, PRE_WORK, \INDEX[2] , \RSHT_BITS[3] , SIGN_Y, C152_DATA4_0,
         C152_DATA4_1, C152_DATA4_2, C152_DATA4_3, C152_DATA4_4, C152_DATA4_5,
         C152_DATA4_6, C152_DATA4_7, C152_DATA4_8, C152_DATA4_9, C152_DATA4_10,
         C152_DATA4_11, N74, N90, N91, N92, N121, N122, N123, N124, N128, N129,
         N657, N658, N659, N660, N661, N662, N663, N664, N665, N666, N667,
         N668, N669, N670, N671, N672, N673, N674, N675, N676, N677, N678,
         N679, N680, N681, N682, N683, N684, N685, N686, N687, N688, N689,
         N690, N691, N692, N693, N694, N695, N696, N697, N698, N699, N700,
         N701, N702, N703, N704, N705, N706, N707, N708, N709, N710, N711,
         N712, N713, N714, N715, N716, N717, N718, N719, N720, N721, N722,
         N723, N724, N725, N726, C2_Z_11, C2_Z_10, C2_Z_9, C2_Z_8, C2_Z_7,
         C2_Z_6, C2_Z_5, C2_Z_4, C2_Z_3, C2_Z_2, C2_Z_1,
         DP_OP_333_124_4748_N57, DP_OP_333_124_4748_N28,
         DP_OP_333_124_4748_N27, DP_OP_333_124_4748_N26,
         DP_OP_333_124_4748_N25, DP_OP_333_124_4748_N24,
         DP_OP_333_124_4748_N23, DP_OP_333_124_4748_N22,
         DP_OP_333_124_4748_N21, DP_OP_333_124_4748_N20,
         DP_OP_333_124_4748_N19, DP_OP_333_124_4748_N18,
         DP_OP_333_124_4748_N12, DP_OP_333_124_4748_N11,
         DP_OP_333_124_4748_N10, DP_OP_333_124_4748_N9, DP_OP_333_124_4748_N8,
         DP_OP_333_124_4748_N7, DP_OP_333_124_4748_N6, DP_OP_333_124_4748_N5,
         DP_OP_333_124_4748_N4, DP_OP_333_124_4748_N3, DP_OP_333_124_4748_N2,
         DP_OP_333_124_4748_N1, INTADD_0_CI, \INTADD_0_SUM[6] ,
         \INTADD_0_SUM[5] , \INTADD_0_SUM[4] , \INTADD_0_SUM[3] ,
         \INTADD_0_SUM[2] , \INTADD_0_SUM[1] , \INTADD_0_SUM[0] , INTADD_0_N7,
         INTADD_0_N6, INTADD_0_N5, INTADD_0_N4, INTADD_0_N3, INTADD_0_N2,
         INTADD_0_N1, ADD_X_132_1_N13, ADD_X_132_1_N12, ADD_X_132_1_N11,
         ADD_X_132_1_N10, ADD_X_132_1_N9, ADD_X_132_1_N8, ADD_X_132_1_N7,
         ADD_X_132_1_N6, ADD_X_132_1_N5, ADD_X_132_1_N4, ADD_X_132_1_N3,
         ADD_X_132_1_N2, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12,
         N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26,
         N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40,
         N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54,
         N55, N56, N57, N58, N59, N60, N61, N63, N103, N104, N105, N106, N107,
         N108, N109, N110, N111, N112, N113, N114, N115, N116, N117, N118,
         N119, N120, N125, N126, N127, N130, N131, N132, N133, N134, N135,
         N136, N137, N138, N139, N140, N141, N142, N143, N144, N145, N146,
         N147, N148, N149, N150, N151, N152, N153, N154, N155, N156, N157,
         N158, N159, N160, N161, N162, N163, N164, N165, N166, N167, N168,
         N169, N170, N171, N172, N173, N174, N175, N176, N177, N178, N179,
         N180, N181, N182, N183, N184, N185, N186, N187, N188, N189, N190,
         N191, N192, N193, N194, N195, N196, N197, N198, N199, N200, N201,
         N202, N203, N204, N205, N206, N207, N208, N209, N210, N211, N212,
         N213, N214, N215, N216, N217, N218, N219, N220, N221, N222, N223,
         N224, N225, N226, N227, N228, N229, N230, N231, N232, N233, N234,
         N235, N236, N237, N238, N239, N240, N241, N242, N243, N244, N245,
         N246, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256,
         N257, N258, N259, N260, N261, N262, N263, N264, N265, N266, N267,
         N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278,
         N279, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289,
         N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300,
         N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311,
         N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322,
         N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333,
         N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344,
         N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355,
         N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, N366,
         N367, N368, N369, N370, N371, N372, N373, N374, N375, N376, N377,
         N378, N379, N380, N381, N382, N383, N384, N385, N386, N387, N388,
         N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399,
         N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410,
         N411, N412, N413, N414, N415, N416, N417, N418, N419, N420, N421,
         N422, N423, N424, N425, N426, N427, N428, N429, N430, N431, N432,
         N433, N434, N435, N436, N437, N438, N439, N440, N441, N442, N443,
         N444, N445, N446, N447, N448, N449, N450, N451, N452, N453, N454,
         N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, N465,
         N466, N467, N468, N469, N470, N471, N472, N473, N474, N475, N476,
         N477, N478, N479, N480, N481, N482, N483, N484, N485, N486, N487,
         N488, N489, N490, N491, N492, N493, N494, N495, N496, N497, N498,
         N499, N500, N501, N502, N503, N504, N505, N506, N507, N508, N509,
         N510, N511, N512, N513, N514, N515, N516, N517, N518, N519, N520,
         N521, N522, N523, N524, N525, N526, N527, N528, N529, N530, N531,
         N532, N533, N534, N535, N536, N537, N538, N539, N540, N541, N542,
         N543, N544, N545, N546, N547, N548, N549, N550, N551, N552, N553,
         N554, N555, N556, N557, N558, N559, N560, N561, N562, N563, N564,
         N565, N566, N567, N568, N569, N570, N571, N572, N573, N574, N575,
         N576, N577, N578, N579, N580, N581, N582, N583, N584, N585, N586,
         N587, N588, N589, N590, N591, N592, N593, N594, N595, N596, N597,
         N598, N599, N600, N601, N602, N603, N604, N605, N606, N607, N608,
         N609, N610, N611, N612, N613, N614, N615, N616, N617, N618, N619,
         N620, N621, N622, N623, N624, N625, N626, N627, N628, N629, N630,
         N631, N632, N633, N634, N635, N636, N637, N638, N639, N640, N641,
         N642, N643, N644, N645, N646, N647, N648, N649, N650, N651, N652,
         N653, N654, N655, N656, N727, N728, N729, N730, N731, N732, N733,
         N734, N735, N736, N737, N738, N739, N740, N741, N742, N743, N744,
         N745, N746, N747, N748, N749, N750, N751, N752, N753, N754, N755,
         N756, N757, N758, N759, N760, N761, N762, N763, N764, N765, N766,
         N767, N768, N769, N770, N771, N772, N773, N774, N775, N776, N777,
         N778, N779, N780, N781, N782, N783, N784, N785, N786, N787, N788,
         N789, N790, N791, N792, N793, N794, N795, N796, N797, N798, N799,
         N800, N801, N802, N803, N804, N805, N806, N807, N808, N809, N810,
         N811, N812, N813, N814, N815, N816, N817, N818, N819, N820, N821,
         N822, N823, N824, N825, N826, N827, N828, N829, N830, N831, N832,
         N833, N834, N835, N836, N837, N838, N839, N840, N841, N842, N843,
         N844, N845, N846, N847, N848, N849, N850, N851, N852, N853, N854,
         N855, N856, N857, N858, N859, N860, N861, N862, N863, N864, N865,
         N866, N867, N868, N869, N870, N871, N872, N873, N874, N875, N876,
         N877, N878, N879, N880, N881, N882, N883, N884, N885, N886, N887,
         N888, N889, N890, N891, N892, N893, N894, N895, N896, N897, N898,
         N899, N900, N901, N902, N903, N904, N905, N906, N907, N908, N909,
         N910, N911, N912, N913, N914, N915, N916, N917, N918, N919, N920,
         N921, N922, N923, N924, N925, N926, N927, N928, N929, N930, N931,
         N932, N933, N934, N935, N936, N937, N938, N939, N940, N941, N942,
         N943, N944, N945, N946, N947, N948, N949, N950, N951, N952, N953,
         N954, N955, N956, N957, N958, N959, N960, N961, N962, N963, N964,
         N965, N966, N967, N968, N969, N970, N971, N972, N973, N974, N975,
         N976, N977, N978, N979, N980, N981, N982, N983, N984, N985, N986,
         N987, N988, N989, N990, N991, N992, N993, N994, N995, N996, N997,
         N998, N999, N1000, N1001, N1002, N1003, N1004, N1005, N1006, N1007,
         N1008, N1009, N1010, N1011, N1012, N1013, N1014, N1015, N1016, N1017,
         N1018, N1019, N1020, N1021, N1022, N1023, N1024, N1025, N1026, N1027,
         N1028, N1029, N1030, N1031, N1032, N1033, N1034, N1035, N1036;
  wire   [12:9] XTEMP;
  wire   [12:0] DIVISION_HEAD;
  wire   [8:0] DIVISION_REMA;
  wire   [12:0] OPER_A;
  wire   [12:0] OPER_B;
  wire   [12:0] SUM_AB;
  wire   [12:0] ZTEMP;
  wire   [3:2] STEP;

  XOR2X1TF \DP_OP_333_124_4748/U27  ( .A(N104), .B(C2_Z_1), .Y(
        DP_OP_333_124_4748_N28) );
  XOR2X1TF \DP_OP_333_124_4748/U26  ( .A(N104), .B(C2_Z_2), .Y(
        DP_OP_333_124_4748_N27) );
  XOR2X1TF \DP_OP_333_124_4748/U25  ( .A(N104), .B(C2_Z_3), .Y(
        DP_OP_333_124_4748_N26) );
  XOR2X1TF \DP_OP_333_124_4748/U24  ( .A(N988), .B(C2_Z_4), .Y(
        DP_OP_333_124_4748_N25) );
  XOR2X1TF \DP_OP_333_124_4748/U23  ( .A(N104), .B(C2_Z_5), .Y(
        DP_OP_333_124_4748_N24) );
  XOR2X1TF \DP_OP_333_124_4748/U22  ( .A(N988), .B(C2_Z_6), .Y(
        DP_OP_333_124_4748_N23) );
  XOR2X1TF \DP_OP_333_124_4748/U21  ( .A(N104), .B(C2_Z_7), .Y(
        DP_OP_333_124_4748_N22) );
  XOR2X1TF \DP_OP_333_124_4748/U20  ( .A(N988), .B(C2_Z_8), .Y(
        DP_OP_333_124_4748_N21) );
  XOR2X1TF \DP_OP_333_124_4748/U19  ( .A(N104), .B(C2_Z_9), .Y(
        DP_OP_333_124_4748_N20) );
  XOR2X1TF \DP_OP_333_124_4748/U18  ( .A(N988), .B(C2_Z_10), .Y(
        DP_OP_333_124_4748_N19) );
  XOR2X1TF \DP_OP_333_124_4748/U17  ( .A(N104), .B(C2_Z_11), .Y(
        DP_OP_333_124_4748_N18) );
  ADDHXLTF \DP_OP_333_124_4748/U12  ( .A(DP_OP_333_124_4748_N28), .B(
        DP_OP_333_124_4748_N12), .CO(DP_OP_333_124_4748_N11), .S(C152_DATA4_1)
         );
  ADDHXLTF \DP_OP_333_124_4748/U11  ( .A(DP_OP_333_124_4748_N27), .B(
        DP_OP_333_124_4748_N11), .CO(DP_OP_333_124_4748_N10), .S(C152_DATA4_2)
         );
  ADDHXLTF \DP_OP_333_124_4748/U10  ( .A(DP_OP_333_124_4748_N26), .B(
        DP_OP_333_124_4748_N10), .CO(DP_OP_333_124_4748_N9), .S(C152_DATA4_3)
         );
  ADDHXLTF \DP_OP_333_124_4748/U9  ( .A(DP_OP_333_124_4748_N25), .B(
        DP_OP_333_124_4748_N9), .CO(DP_OP_333_124_4748_N8), .S(C152_DATA4_4)
         );
  ADDHXLTF \DP_OP_333_124_4748/U8  ( .A(DP_OP_333_124_4748_N24), .B(
        DP_OP_333_124_4748_N8), .CO(DP_OP_333_124_4748_N7), .S(C152_DATA4_5)
         );
  ADDHXLTF \DP_OP_333_124_4748/U7  ( .A(DP_OP_333_124_4748_N23), .B(
        DP_OP_333_124_4748_N7), .CO(DP_OP_333_124_4748_N6), .S(C152_DATA4_6)
         );
  ADDHXLTF \DP_OP_333_124_4748/U6  ( .A(DP_OP_333_124_4748_N22), .B(
        DP_OP_333_124_4748_N6), .CO(DP_OP_333_124_4748_N5), .S(C152_DATA4_7)
         );
  ADDHXLTF \DP_OP_333_124_4748/U5  ( .A(DP_OP_333_124_4748_N21), .B(
        DP_OP_333_124_4748_N5), .CO(DP_OP_333_124_4748_N4), .S(C152_DATA4_8)
         );
  ADDHXLTF \DP_OP_333_124_4748/U4  ( .A(DP_OP_333_124_4748_N20), .B(
        DP_OP_333_124_4748_N4), .CO(DP_OP_333_124_4748_N3), .S(C152_DATA4_9)
         );
  ADDHXLTF \DP_OP_333_124_4748/U3  ( .A(DP_OP_333_124_4748_N19), .B(
        DP_OP_333_124_4748_N3), .CO(DP_OP_333_124_4748_N2), .S(C152_DATA4_10)
         );
  ADDHXLTF \DP_OP_333_124_4748/U2  ( .A(DP_OP_333_124_4748_N18), .B(
        DP_OP_333_124_4748_N2), .CO(DP_OP_333_124_4748_N1), .S(C152_DATA4_11)
         );
  CMPR32X2TF \intadd_0/U8  ( .A(X_IN[1]), .B(DIVISION_HEAD[5]), .C(INTADD_0_CI), .CO(INTADD_0_N7), .S(\INTADD_0_SUM[0] ) );
  CMPR32X2TF \intadd_0/U7  ( .A(X_IN[2]), .B(DIVISION_HEAD[6]), .C(INTADD_0_N7), .CO(INTADD_0_N6), .S(\INTADD_0_SUM[1] ) );
  CMPR32X2TF \intadd_0/U6  ( .A(X_IN[3]), .B(DIVISION_HEAD[7]), .C(INTADD_0_N6), .CO(INTADD_0_N5), .S(\INTADD_0_SUM[2] ) );
  CMPR32X2TF \intadd_0/U5  ( .A(X_IN[4]), .B(DIVISION_HEAD[8]), .C(INTADD_0_N5), .CO(INTADD_0_N4), .S(\INTADD_0_SUM[3] ) );
  CMPR32X2TF \intadd_0/U4  ( .A(X_IN[5]), .B(DIVISION_HEAD[9]), .C(INTADD_0_N4), .CO(INTADD_0_N3), .S(\INTADD_0_SUM[4] ) );
  CMPR32X2TF \intadd_0/U3  ( .A(X_IN[6]), .B(DIVISION_HEAD[10]), .C(
        INTADD_0_N3), .CO(INTADD_0_N2), .S(\INTADD_0_SUM[5] ) );
  CMPR32X2TF \intadd_0/U2  ( .A(X_IN[7]), .B(DIVISION_HEAD[11]), .C(
        INTADD_0_N2), .CO(INTADD_0_N1), .S(\INTADD_0_SUM[6] ) );
  DFFRX2TF \wtemp_reg[9]  ( .D(N673), .CK(CLK), .RN(RST_N), .Q(OPER_B[9]), 
        .QN(N202) );
  DFFRX2TF \wtemp_reg[12]  ( .D(N724), .CK(CLK), .RN(RST_N), .Q(OPER_B[12]), 
        .QN(N201) );
  DFFRX2TF \wtemp_reg[11]  ( .D(N671), .CK(CLK), .RN(RST_N), .Q(OPER_B[11]), 
        .QN(N199) );
  DFFRX2TF \wtemp_reg[0]  ( .D(N682), .CK(CLK), .RN(RST_N), .Q(OPER_B[0]), 
        .QN(N198) );
  DFFRX2TF \wtemp_reg[3]  ( .D(N679), .CK(CLK), .RN(RST_N), .Q(OPER_B[3]), 
        .QN(N197) );
  DFFRX2TF \wtemp_reg[1]  ( .D(N681), .CK(CLK), .RN(RST_N), .Q(OPER_B[1]), 
        .QN(N196) );
  DFFRX2TF \wtemp_reg[4]  ( .D(N678), .CK(CLK), .RN(RST_N), .Q(OPER_B[4]), 
        .QN(N191) );
  DFFSX2TF pre_work_reg ( .D(N695), .CK(CLK), .SN(RST_N), .Q(PRE_WORK), .QN(
        N190) );
  DFFRX2TF \ytemp_reg[1]  ( .D(N693), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[1]), .QN(N184) );
  DFFRX2TF \ytemp_reg[2]  ( .D(N692), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[2]), .QN(N180) );
  DFFRX2TF \xtemp_reg[0]  ( .D(N719), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[4]), .QN(N179) );
  DFFRX2TF \xtemp_reg[10]  ( .D(N709), .CK(CLK), .RN(RST_N), .Q(XTEMP[10]), 
        .QN(N176) );
  DFFRX2TF \xtemp_reg[8]  ( .D(N711), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[12]), .QN(N175) );
  DFFRX2TF \ytemp_reg[6]  ( .D(N688), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[6]), .QN(N174) );
  DFFRX2TF \ytemp_reg[4]  ( .D(N690), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[4]), .QN(N173) );
  DFFRX2TF \ytemp_reg[9]  ( .D(N685), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[0]), .QN(N172) );
  DFFRX2TF \ytemp_reg[7]  ( .D(N687), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[7]), .QN(N171) );
  DFFRX2TF \ytemp_reg[5]  ( .D(N689), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[5]), .QN(N170) );
  DFFRX2TF \xtemp_reg[11]  ( .D(N708), .CK(CLK), .RN(RST_N), .Q(XTEMP[11]), 
        .QN(N169) );
  DFFRX2TF \xtemp_reg[3]  ( .D(N716), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[7]), .QN(N168) );
  DFFRX2TF \xtemp_reg[2]  ( .D(N717), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[6]), .QN(N167) );
  DFFRX2TF \ytemp_reg[10]  ( .D(N684), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[1]), .QN(N165) );
  DFFRX2TF \ytemp_reg[8]  ( .D(N686), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[8]), .QN(N164) );
  ADDHX1TF \add_x_132_1/U14  ( .A(OPER_B[0]), .B(OPER_A[0]), .CO(
        ADD_X_132_1_N13), .S(SUM_AB[0]) );
  CMPR32X2TF \add_x_132_1/U4  ( .A(OPER_A[10]), .B(OPER_B[10]), .C(
        ADD_X_132_1_N4), .CO(ADD_X_132_1_N3), .S(SUM_AB[10]) );
  CMPR32X2TF \add_x_132_1/U6  ( .A(OPER_A[8]), .B(OPER_B[8]), .C(
        ADD_X_132_1_N6), .CO(ADD_X_132_1_N5), .S(SUM_AB[8]) );
  CMPR32X2TF \add_x_132_1/U10  ( .A(OPER_A[4]), .B(OPER_B[4]), .C(
        ADD_X_132_1_N10), .CO(ADD_X_132_1_N9), .S(SUM_AB[4]) );
  CMPR32X2TF \add_x_132_1/U12  ( .A(OPER_A[2]), .B(OPER_B[2]), .C(
        ADD_X_132_1_N12), .CO(ADD_X_132_1_N11), .S(SUM_AB[2]) );
  CMPR32X2TF \add_x_132_1/U13  ( .A(OPER_A[1]), .B(OPER_B[1]), .C(
        ADD_X_132_1_N13), .CO(ADD_X_132_1_N12), .S(SUM_AB[1]) );
  CMPR32X2TF \add_x_132_1/U5  ( .A(OPER_A[9]), .B(OPER_B[9]), .C(
        ADD_X_132_1_N5), .CO(ADD_X_132_1_N4), .S(SUM_AB[9]) );
  CMPR32X2TF \add_x_132_1/U11  ( .A(OPER_A[3]), .B(OPER_B[3]), .C(
        ADD_X_132_1_N11), .CO(ADD_X_132_1_N10), .S(SUM_AB[3]) );
  CMPR32X2TF \add_x_132_1/U9  ( .A(OPER_A[5]), .B(OPER_B[5]), .C(
        ADD_X_132_1_N9), .CO(ADD_X_132_1_N8), .S(SUM_AB[5]) );
  CMPR32X2TF \add_x_132_1/U3  ( .A(OPER_A[11]), .B(OPER_B[11]), .C(
        ADD_X_132_1_N3), .CO(ADD_X_132_1_N2), .S(SUM_AB[11]) );
  DFFRX1TF \rsht_bits_reg[2]  ( .D(N701), .CK(CLK), .RN(RST_N), .QN(N90) );
  DFFSRX2TF sign_y_reg ( .D(N694), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(SIGN_Y), 
        .QN(N192) );
  DFFSRX2TF XOR_SRC_reg ( .D(N707), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(N61), 
        .QN(N130) );
  DFFSRX2TF \rsht_bits_reg[0]  ( .D(N703), .CK(CLK), .SN(1'b1), .RN(RST_N), 
        .Q(N194), .QN(N92) );
  DFFSRX2TF \step_reg[1]  ( .D(N700), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(N177), .QN(N121) );
  DFFSRX2TF \step_reg[3]  ( .D(N721), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        STEP[3]), .QN(N178) );
  DFFSRX2TF \step_reg[2]  ( .D(N696), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        STEP[2]), .QN(N166) );
  DFFSRX2TF \rsht_bits_reg[1]  ( .D(N702), .CK(CLK), .SN(1'b1), .RN(RST_N), 
        .Q(N183), .QN(N91) );
  DFFSRX2TF \step_reg[0]  ( .D(N697), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(N188), .QN(N122) );
  DFFSRX2TF \rsht_bits_reg[3]  ( .D(N704), .CK(CLK), .SN(1'b1), .RN(RST_N), 
        .Q(\RSHT_BITS[3] ), .QN(N203) );
  DFFSRX2TF SEL_SRC_reg ( .D(N720), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        POST_WORK), .QN(N187) );
  DFFSRX2TF \index_reg[1]  ( .D(N699), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        N195), .QN(N128) );
  DFFSRX2TF SEL_Z_reg ( .D(N670), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(N189), 
        .QN(N123) );
  DFFSRX2TF \index_reg[3]  ( .D(N725), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        N200), .QN(N124) );
  DFFSRX2TF \index_reg[0]  ( .D(N726), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        N182), .QN(N129) );
  DFFSRX2TF \ytemp_reg[0]  ( .D(N705), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        DIVISION_REMA[0]), .QN(N193) );
  DFFSRX2TF \wtemp_reg[8]  ( .D(N674), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        OPER_B[8]), .QN(N185) );
  DFFSRX2TF \wtemp_reg[2]  ( .D(N680), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        OPER_B[2]), .QN(N181) );
  DFFSRX2TF \wtemp_reg[10]  ( .D(N672), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        OPER_B[10]), .QN(N186) );
  DFFRX1TF \ztemp_reg[0]  ( .D(N669), .CK(CLK), .RN(RST_N), .Q(ZTEMP[0]) );
  DFFRX1TF \wtemp_reg[6]  ( .D(N676), .CK(CLK), .RN(RST_N), .Q(OPER_B[6]) );
  DFFRX1TF \ztemp_reg[8]  ( .D(N661), .CK(CLK), .RN(RST_N), .Q(ZTEMP[8]) );
  DFFRX1TF \ztemp_reg[6]  ( .D(N663), .CK(CLK), .RN(RST_N), .Q(ZTEMP[6]) );
  DFFRX1TF \ztemp_reg[4]  ( .D(N665), .CK(CLK), .RN(RST_N), .Q(ZTEMP[4]) );
  DFFRX1TF \ztemp_reg[2]  ( .D(N667), .CK(CLK), .RN(RST_N), .Q(ZTEMP[2]) );
  DFFRX1TF \ztemp_reg[1]  ( .D(N668), .CK(CLK), .RN(RST_N), .Q(ZTEMP[1]) );
  DFFRX1TF \ztemp_reg[5]  ( .D(N664), .CK(CLK), .RN(RST_N), .Q(ZTEMP[5]) );
  DFFRX1TF \ztemp_reg[3]  ( .D(N666), .CK(CLK), .RN(RST_N), .Q(ZTEMP[3]) );
  DFFRX1TF \ztemp_reg[7]  ( .D(N662), .CK(CLK), .RN(RST_N), .Q(ZTEMP[7]) );
  DFFRX1TF \ztemp_reg[9]  ( .D(N660), .CK(CLK), .RN(RST_N), .Q(ZTEMP[9]) );
  DFFRX1TF \ytemp_reg[3]  ( .D(N691), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[3]), .QN(N752) );
  DFFRX1TF \wtemp_reg[5]  ( .D(N677), .CK(CLK), .RN(RST_N), .Q(OPER_B[5]) );
  DFFRX1TF \wtemp_reg[7]  ( .D(N675), .CK(CLK), .RN(RST_N), .Q(OPER_B[7]) );
  DFFRX1TF \ztemp_reg[10]  ( .D(N659), .CK(CLK), .RN(RST_N), .Q(ZTEMP[10]) );
  DFFRX1TF \ztemp_reg[11]  ( .D(N658), .CK(CLK), .RN(RST_N), .Q(ZTEMP[11]) );
  DFFRX1TF \ztemp_reg[12]  ( .D(N657), .CK(CLK), .RN(RST_N), .Q(ZTEMP[12]) );
  DFFRX1TF \xtemp_reg[12]  ( .D(N723), .CK(CLK), .RN(RST_N), .Q(XTEMP[12]), 
        .QN(N368) );
  DFFRX1TF \ytemp_reg[11]  ( .D(N683), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[2]), .QN(N829) );
  DFFRX1TF \ytemp_reg[12]  ( .D(N706), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[3]), .QN(N734) );
  DFFRX2TF \xtemp_reg[1]  ( .D(N718), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[5]), .QN(N527) );
  DFFRX2TF \xtemp_reg[9]  ( .D(N710), .CK(CLK), .RN(RST_N), .Q(XTEMP[9]), .QN(
        N544) );
  DFFRX2TF \xtemp_reg[7]  ( .D(N712), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[11]), .QN(N477) );
  DFFRX2TF \xtemp_reg[5]  ( .D(N714), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[9]), .QN(N455) );
  DFFRX2TF \xtemp_reg[6]  ( .D(N713), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[10]), .QN(N541) );
  DFFRX2TF \xtemp_reg[4]  ( .D(N715), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[8]), .QN(N536) );
  DFFRX2TF sign_x_reg ( .D(N722), .CK(CLK), .RN(RST_N), .Q(N982), .QN(N74) );
  DFFRX2TF \index_reg[2]  ( .D(N698), .CK(CLK), .RN(RST_N), .Q(\INDEX[2] ) );
  OA21XLTF U3 ( .A0(SUM_AB[12]), .A1(N736), .B0(N145), .Y(N160) );
  NAND2X1TF U4 ( .A(PRE_WORK), .B(N988), .Y(N398) );
  CLKBUFX2TF U5 ( .A(N271), .Y(N204) );
  CLKBUFX2TF U6 ( .A(N204), .Y(N159) );
  AOI32XLTF U7 ( .A0(N838), .A1(N103), .A2(N839), .B0(N653), .B1(N958), .Y(
        N729) );
  AOI211X2TF U8 ( .A0(N586), .A1(N103), .B0(N610), .C0(N585), .Y(N612) );
  AND2X2TF U9 ( .A(N231), .B(PRE_WORK), .Y(DP_OP_333_124_4748_N57) );
  AOI21X1TF U10 ( .A0(N842), .A1(N948), .B0(N865), .Y(N1) );
  NOR3X1TF U11 ( .A(OPER_A[1]), .B(N951), .C(N842), .Y(N2) );
  OAI32X1TF U12 ( .A0(N196), .A1(OPER_B[0]), .A2(N141), .B0(N952), .B1(N196), 
        .Y(N3) );
  AOI211X1TF U13 ( .A0(OPER_B[2]), .A1(N875), .B0(N2), .C0(N3), .Y(N4) );
  OAI31X1TF U14 ( .A0(N141), .A1(N198), .A2(OPER_B[1]), .B0(N841), .Y(N5) );
  AOI211X1TF U15 ( .A0(C152_DATA4_1), .A1(N139), .B0(N903), .C0(N5), .Y(N6) );
  OAI211X1TF U16 ( .A0(N843), .A1(N1), .B0(N4), .C0(N6), .Y(N681) );
  AOI22X1TF U17 ( .A0(DIVISION_HEAD[0]), .A1(N132), .B0(ZTEMP[0]), .B1(N1028), 
        .Y(N7) );
  AOI32XLTF U18 ( .A0(N1036), .A1(N7), .A2(N1027), .B0(N993), .B1(N7), .Y(N669) );
  AOI32X1TF U19 ( .A0(N141), .A1(N854), .A2(N952), .B0(N198), .B1(N854), .Y(N8) );
  AOI211X1TF U20 ( .A0(C152_DATA4_0), .A1(N139), .B0(N903), .C0(N8), .Y(N9) );
  OAI21X1TF U21 ( .A0(N865), .A1(N948), .B0(OPER_A[0]), .Y(N10) );
  OAI211X1TF U22 ( .A0(N196), .A1(N911), .B0(N9), .C0(N10), .Y(N682) );
  NOR3X1TF U23 ( .A(Y_IN[12]), .B(Y_IN[11]), .C(Y_IN[10]), .Y(N11) );
  CLKINVX1TF U24 ( .A(N454), .Y(N12) );
  AOI22X1TF U25 ( .A0(N325), .A1(N12), .B0(N127), .B1(N754), .Y(N13) );
  OAI21X1TF U26 ( .A0(X_IN[4]), .A1(N324), .B0(N114), .Y(N14) );
  OAI22X1TF U27 ( .A0(N127), .A1(N754), .B0(X_IN[6]), .B1(N746), .Y(N15) );
  AOI31X1TF U28 ( .A0(N326), .A1(N13), .A2(N14), .B0(N15), .Y(N16) );
  AOI21X1TF U29 ( .A0(N746), .A1(X_IN[6]), .B0(N16), .Y(N17) );
  OA22X1TF U30 ( .A0(N18), .A1(N17), .B0(N502), .B1(N206), .Y(N19) );
  AO21X1TF U31 ( .A0(N482), .A1(N17), .B0(Y_IN[4]), .Y(N20) );
  AOI22X1TF U32 ( .A0(N502), .A1(N206), .B0(N19), .B1(N20), .Y(N21) );
  AOI2BB2X1TF U33 ( .B0(X_IN[9]), .B1(N21), .A0N(N515), .A1N(N113), .Y(N22) );
  CLKINVX1TF U34 ( .A(N21), .Y(N23) );
  AO21X1TF U35 ( .A0(N514), .A1(N23), .B0(Y_IN[6]), .Y(N24) );
  AOI22X1TF U36 ( .A0(N515), .A1(N113), .B0(N22), .B1(N24), .Y(N25) );
  AOI222XLTF U37 ( .A0(N778), .A1(X_IN[11]), .B0(N778), .B1(N25), .C0(X_IN[11]), .C1(N25), .Y(N26) );
  OAI21X1TF U38 ( .A0(Y_IN[9]), .A1(N315), .B0(N26), .Y(N27) );
  OAI211X1TF U39 ( .A0(X_IN[12]), .A1(N800), .B0(N11), .C0(N27), .Y(N786) );
  CLKINVX1TF U40 ( .A(X_IN[7]), .Y(N18) );
  OAI32X1TF U41 ( .A0(N199), .A1(N953), .A2(N141), .B0(N952), .B1(N199), .Y(
        N28) );
  CLKINVX1TF U42 ( .A(OPER_A[11]), .Y(N29) );
  OAI32X1TF U43 ( .A0(N29), .A1(N951), .A2(N950), .B0(N949), .B1(N29), .Y(N30)
         );
  AOI31X1TF U44 ( .A0(N950), .A1(N948), .A2(N29), .B0(N947), .Y(N31) );
  NOR2X1TF U45 ( .A(N140), .B(OPER_B[11]), .Y(N32) );
  AOI222XLTF U46 ( .A0(C152_DATA4_11), .A1(N138), .B0(N233), .B1(N981), .C0(
        N953), .C1(N32), .Y(N33) );
  OAI211X1TF U47 ( .A0(N201), .A1(N955), .B0(N31), .C0(N33), .Y(N34) );
  OR3X1TF U48 ( .A(N28), .B(N30), .C(N34), .Y(N671) );
  OAI21X1TF U49 ( .A0(N322), .A1(N644), .B0(N637), .Y(N35) );
  AND4X1TF U50 ( .A(\INDEX[2] ), .B(N640), .C(N633), .D(N124), .Y(N36) );
  AOI211X1TF U51 ( .A0(N200), .A1(N35), .B0(N36), .C0(N394), .Y(N37) );
  NAND3X1TF U52 ( .A(N372), .B(N820), .C(N37), .Y(N725) );
  NOR2X1TF U53 ( .A(N950), .B(OPER_A[11]), .Y(N38) );
  XNOR2X1TF U54 ( .A(OPER_A[12]), .B(N38), .Y(N39) );
  AOI22X1TF U55 ( .A0(N39), .A1(N948), .B0(OPER_A[12]), .B1(N865), .Y(N40) );
  OAI21X1TF U56 ( .A0(N152), .A1(N564), .B0(N143), .Y(N41) );
  XNOR2X1TF U57 ( .A(N41), .B(N104), .Y(N42) );
  XNOR2X1TF U58 ( .A(DP_OP_333_124_4748_N1), .B(N42), .Y(N43) );
  NOR2X1TF U59 ( .A(OPER_B[11]), .B(N953), .Y(N44) );
  OAI31X1TF U60 ( .A0(N140), .A1(N44), .A2(OPER_B[12]), .B0(N841), .Y(N45) );
  AOI211X1TF U61 ( .A0(N139), .A1(N43), .B0(N947), .C0(N45), .Y(N46) );
  OAI31X1TF U62 ( .A0(OPER_B[11]), .A1(N953), .A2(N928), .B0(N885), .Y(N47) );
  AOI32X1TF U63 ( .A0(N958), .A1(OPER_B[12]), .A2(N47), .B0(N230), .B1(
        OPER_B[12]), .Y(N48) );
  NAND4BX1TF U64 ( .AN(N837), .B(N40), .C(N46), .D(N48), .Y(N724) );
  OAI21X1TF U65 ( .A0(N151), .A1(N742), .B0(N142), .Y(N49) );
  CLKMX2X2TF U66 ( .A(N104), .B(DP_OP_333_124_4748_N57), .S0(N49), .Y(
        DP_OP_333_124_4748_N12) );
  XOR2X1TF U67 ( .A(DP_OP_333_124_4748_N57), .B(N49), .Y(C152_DATA4_0) );
  NOR3X1TF U68 ( .A(N927), .B(N74), .C(N924), .Y(N50) );
  NOR2X1TF U69 ( .A(N186), .B(N955), .Y(N51) );
  AOI211X1TF U70 ( .A0(N138), .A1(C152_DATA4_9), .B0(N50), .C0(N51), .Y(N52)
         );
  NOR2X1TF U71 ( .A(N951), .B(OPER_A[9]), .Y(N53) );
  AOI22X1TF U72 ( .A0(SIGN_Y), .A1(N923), .B0(N926), .B1(N53), .Y(N54) );
  OAI21X1TF U73 ( .A0(N141), .A1(N925), .B0(N952), .Y(N55) );
  OAI21X1TF U74 ( .A0(N951), .A1(N926), .B0(N949), .Y(N56) );
  AOI22X1TF U75 ( .A0(OPER_B[9]), .A1(N55), .B0(OPER_A[9]), .B1(N56), .Y(N57)
         );
  NAND3X1TF U76 ( .A(N954), .B(N925), .C(N202), .Y(N58) );
  NAND4X1TF U77 ( .A(N52), .B(N54), .C(N57), .D(N58), .Y(N673) );
  OR2X2TF U78 ( .A(N358), .B(N615), .Y(N59) );
  INVX2TF U79 ( .A(N988), .Y(N151) );
  INVX2TF U80 ( .A(N958), .Y(N144) );
  INVX2TF U81 ( .A(N144), .Y(N103) );
  OR3X1TF U82 ( .A(PRE_WORK), .B(N621), .C(N615), .Y(N60) );
  NAND2X2TF U83 ( .A(SIGN_Y), .B(N982), .Y(N989) );
  AOI22XLTF U84 ( .A0(DIVISION_HEAD[10]), .A1(N563), .B0(DIVISION_HEAD[9]), 
        .B1(N800), .Y(N339) );
  INVX2TF U85 ( .A(N123), .Y(N63) );
  NAND2X1TF U104 ( .A(N790), .B(N782), .Y(N407) );
  NAND2X1TF U105 ( .A(N946), .B(N215), .Y(N229) );
  NAND2XLTF U106 ( .A(N816), .B(SUM_AB[8]), .Y(N436) );
  CLKINVX1TF U107 ( .A(SUM_AB[4]), .Y(N401) );
  AO21X1TF U108 ( .A0(N793), .A1(N384), .B0(N839), .Y(N522) );
  CLKINVX2TF U109 ( .A(OPER_A[4]), .Y(N873) );
  CLKINVX1TF U110 ( .A(N878), .Y(N876) );
  AND2X2TF U111 ( .A(ZTEMP[5]), .B(N204), .Y(POUT[5]) );
  AND2X2TF U112 ( .A(ZTEMP[6]), .B(N204), .Y(POUT[6]) );
  CLKINVX1TF U113 ( .A(N850), .Y(N845) );
  CLKINVX1TF U114 ( .A(N636), .Y(N638) );
  CLKINVX1TF U115 ( .A(N206), .Y(N213) );
  CLKBUFX2TF U116 ( .A(ALU_START), .Y(N106) );
  CLKINVX1TF U117 ( .A(Y_IN[6]), .Y(N212) );
  CLKINVX1TF U118 ( .A(X_IN[2]), .Y(N788) );
  AOI211X1TF U119 ( .A0(X_IN[3]), .A1(N763), .B0(N452), .C0(N451), .Y(N453) );
  AOI211X1TF U120 ( .A0(X_IN[5]), .A1(N763), .B0(N471), .C0(N470), .Y(N472) );
  AOI211X1TF U121 ( .A0(Y_IN[7]), .A1(N763), .B0(N804), .C0(N803), .Y(N805) );
  OA21XLTF U122 ( .A0(SUM_AB[12]), .A1(N406), .B0(N145), .Y(N518) );
  CLKINVX2TF U123 ( .A(N882), .Y(N223) );
  INVX1TF U124 ( .A(N923), .Y(N900) );
  AND2X2TF U125 ( .A(N921), .B(N939), .Y(N954) );
  OR2X2TF U126 ( .A(N1028), .B(N151), .Y(N1029) );
  OAI31X1TF U127 ( .A0(N295), .A1(X_IN[11]), .A2(N563), .B0(N294), .Y(N296) );
  AOI22X1TF U128 ( .A0(X_IN[5]), .A1(N457), .B0(N105), .B1(N125), .Y(N459) );
  AOI22X1TF U129 ( .A0(Y_IN[9]), .A1(N818), .B0(X_IN[4]), .B1(N155), .Y(N819)
         );
  AOI22X1TF U130 ( .A0(X_IN[2]), .A1(N155), .B0(X_IN[3]), .B1(N823), .Y(N802)
         );
  AOI22X1TF U131 ( .A0(X_IN[12]), .A1(N823), .B0(X_IN[11]), .B1(N155), .Y(N448) );
  OAI21X1TF U132 ( .A0(N390), .A1(N763), .B0(N392), .Y(N391) );
  AOI22X1TF U133 ( .A0(XTEMP[11]), .A1(N150), .B0(N105), .B1(N457), .Y(N364)
         );
  AOI21X1TF U134 ( .A0(N728), .A1(N958), .B0(N727), .Y(N731) );
  INVX1TF U135 ( .A(N416), .Y(N417) );
  NAND3XLTF U136 ( .A(N958), .B(N840), .C(N839), .Y(N648) );
  OAI31X1TF U137 ( .A0(N580), .A1(N581), .A2(N579), .B0(N103), .Y(N597) );
  NAND4XLTF U138 ( .A(N627), .B(N626), .C(N625), .D(N624), .Y(N628) );
  OR2X2TF U139 ( .A(N398), .B(N780), .Y(N817) );
  OAI2BB2XLTF U140 ( .B0(N778), .B1(N820), .A0N(Y_IN[6]), .A1N(N818), .Y(N795)
         );
  OAI31XLTF U141 ( .A0(N145), .A1(N188), .A2(N647), .B0(N646), .Y(N652) );
  AOI22X1TF U142 ( .A0(Y_IN[1]), .A1(N818), .B0(DIVISION_REMA[4]), .B1(N147), 
        .Y(N747) );
  NAND3BXLTF U143 ( .AN(N393), .B(N793), .C(N654), .Y(N377) );
  OAI211XLTF U144 ( .A0(N152), .A1(N376), .B0(N990), .C0(N616), .Y(N378) );
  AOI22X1TF U145 ( .A0(DIVISION_HEAD[2]), .A1(N147), .B0(Y_IN[8]), .B1(N818), 
        .Y(N811) );
  AOI22X1TF U146 ( .A0(Y_IN[3]), .A1(N818), .B0(DIVISION_REMA[6]), .B1(N147), 
        .Y(N758) );
  AOI22X1TF U147 ( .A0(N206), .A1(N818), .B0(Y_IN[7]), .B1(N807), .Y(N771) );
  AOI22X1TF U148 ( .A0(X_IN[2]), .A1(N457), .B0(X_IN[1]), .B1(N818), .Y(N430)
         );
  INVX1TF U149 ( .A(OPER_A[10]), .Y(N932) );
  INVX1TF U150 ( .A(OPER_A[6]), .Y(N892) );
  INVX1TF U151 ( .A(OPER_A[8]), .Y(N914) );
  INVX2TF U152 ( .A(N751), .Y(N119) );
  INVX1TF U153 ( .A(OPER_A[1]), .Y(N843) );
  INVX2TF U154 ( .A(N763), .Y(N117) );
  INVX2TF U155 ( .A(N151), .Y(N104) );
  AOI22X1TF U156 ( .A0(DIVISION_HEAD[2]), .A1(N135), .B0(ZTEMP[11]), .B1(N63), 
        .Y(N267) );
  AOI22X1TF U157 ( .A0(DIVISION_HEAD[0]), .A1(N135), .B0(ZTEMP[9]), .B1(N63), 
        .Y(N265) );
  AOI22X1TF U158 ( .A0(DIVISION_REMA[8]), .A1(N135), .B0(ZTEMP[8]), .B1(N189), 
        .Y(N264) );
  AOI22X1TF U159 ( .A0(DIVISION_HEAD[1]), .A1(N135), .B0(ZTEMP[10]), .B1(N63), 
        .Y(N266) );
  AOI22X1TF U160 ( .A0(DIVISION_REMA[7]), .A1(N135), .B0(ZTEMP[7]), .B1(N189), 
        .Y(N263) );
  AOI22X1TF U161 ( .A0(DIVISION_REMA[6]), .A1(N135), .B0(ZTEMP[6]), .B1(N189), 
        .Y(N262) );
  AOI22X1TF U162 ( .A0(DIVISION_REMA[5]), .A1(N135), .B0(ZTEMP[5]), .B1(N189), 
        .Y(N261) );
  AOI22X1TF U163 ( .A0(DIVISION_REMA[4]), .A1(N135), .B0(ZTEMP[4]), .B1(N189), 
        .Y(N260) );
  AOI22X1TF U164 ( .A0(DIVISION_REMA[3]), .A1(N135), .B0(ZTEMP[3]), .B1(N189), 
        .Y(N259) );
  AOI22X1TF U165 ( .A0(DIVISION_REMA[2]), .A1(N134), .B0(ZTEMP[2]), .B1(N189), 
        .Y(N258) );
  AOI22X1TF U166 ( .A0(DIVISION_REMA[1]), .A1(N134), .B0(ZTEMP[1]), .B1(N189), 
        .Y(N257) );
  AOI22X1TF U167 ( .A0(DIVISION_REMA[0]), .A1(N134), .B0(ZTEMP[0]), .B1(N189), 
        .Y(N256) );
  CLKAND2X2TF U168 ( .A(N732), .B(N655), .Y(N561) );
  INVX2TF U169 ( .A(N59), .Y(N146) );
  AOI22X1TF U170 ( .A0(DIVISION_HEAD[3]), .A1(N135), .B0(ZTEMP[12]), .B1(N63), 
        .Y(N269) );
  AND2X2TF U171 ( .A(N395), .B(N361), .Y(N751) );
  INVX2TF U172 ( .A(N268), .Y(N134) );
  INVX1TF U173 ( .A(N352), .Y(N972) );
  AND2X2TF U174 ( .A(N352), .B(N231), .Y(N958) );
  AND2X2TF U175 ( .A(N361), .B(DP_OP_333_124_4748_N57), .Y(N763) );
  NAND2XLTF U176 ( .A(N231), .B(N963), .Y(N549) );
  INVX2TF U177 ( .A(N356), .Y(N357) );
  AND2X2TF U178 ( .A(N123), .B(N255), .Y(N270) );
  OR2X2TF U179 ( .A(N189), .B(N255), .Y(N268) );
  INVX2TF U180 ( .A(N207), .Y(N113) );
  AND2X2TF U181 ( .A(N61), .B(N204), .Y(N253) );
  AND2X2TF U182 ( .A(N232), .B(N106), .Y(N988) );
  AND2X2TF U183 ( .A(N204), .B(N130), .Y(N252) );
  INVX2TF U184 ( .A(N209), .Y(N127) );
  AOI22X1TF U185 ( .A0(X_IN[11]), .A1(N563), .B0(X_IN[12]), .B1(N821), .Y(N290) );
  INVX1TF U186 ( .A(N272), .Y(N157) );
  NAND2XLTF U187 ( .A(DIVISION_HEAD[4]), .B(N272), .Y(N234) );
  INVX2TF U188 ( .A(X_IN[3]), .Y(N208) );
  INVX2TF U189 ( .A(X_IN[5]), .Y(N209) );
  INVX2TF U190 ( .A(Y_IN[7]), .Y(N207) );
  INVX2TF U191 ( .A(N311), .Y(N105) );
  INVX2TF U192 ( .A(N253), .Y(N107) );
  INVX2TF U193 ( .A(N253), .Y(N108) );
  INVX2TF U194 ( .A(N252), .Y(N109) );
  INVX2TF U195 ( .A(N252), .Y(N110) );
  INVX2TF U196 ( .A(N1036), .Y(N111) );
  INVX2TF U197 ( .A(N1036), .Y(N112) );
  INVX2TF U198 ( .A(N208), .Y(N114) );
  INVX2TF U199 ( .A(N60), .Y(N115) );
  INVX2TF U200 ( .A(N60), .Y(N116) );
  INVX2TF U201 ( .A(N763), .Y(N118) );
  INVX2TF U202 ( .A(N751), .Y(N120) );
  INVX2TF U203 ( .A(N407), .Y(N125) );
  INVX2TF U204 ( .A(N407), .Y(N126) );
  INVX2TF U205 ( .A(N130), .Y(N131) );
  INVX2TF U206 ( .A(N1029), .Y(N132) );
  INVX2TF U207 ( .A(N1029), .Y(N133) );
  INVX2TF U208 ( .A(N268), .Y(N135) );
  INVX2TF U209 ( .A(N270), .Y(N136) );
  INVX2TF U210 ( .A(N270), .Y(N137) );
  INVX2TF U211 ( .A(N229), .Y(N138) );
  INVX2TF U212 ( .A(N229), .Y(N139) );
  INVX2TF U213 ( .A(N954), .Y(N140) );
  INVX2TF U214 ( .A(N954), .Y(N141) );
  INVX2TF U215 ( .A(DP_OP_333_124_4748_N57), .Y(N142) );
  INVX2TF U216 ( .A(DP_OP_333_124_4748_N57), .Y(N143) );
  INVX2TF U217 ( .A(N958), .Y(N145) );
  INVX2TF U218 ( .A(N59), .Y(N147) );
  INVX2TF U219 ( .A(N522), .Y(N148) );
  INVX2TF U220 ( .A(N522), .Y(N149) );
  INVX2TF U221 ( .A(N119), .Y(N150) );
  INVX2TF U222 ( .A(N988), .Y(N152) );
  AOI222X4TF U223 ( .A0(N501), .A1(N176), .B0(N501), .B1(N515), .C0(N176), 
        .C1(N515), .Y(N511) );
  NOR2X2TF U224 ( .A(N349), .B(N973), .Y(N361) );
  NOR2X2TF U225 ( .A(N358), .B(N151), .Y(N395) );
  NOR3X2TF U226 ( .A(N144), .B(N620), .C(N647), .Y(N633) );
  INVX2TF U227 ( .A(N518), .Y(N153) );
  INVX2TF U228 ( .A(N518), .Y(N154) );
  INVX2TF U229 ( .A(N817), .Y(N155) );
  INVX2TF U230 ( .A(N817), .Y(N156) );
  NAND2X2TF U231 ( .A(N123), .B(N779), .Y(N467) );
  AOI21X2TF U232 ( .A0(N103), .A1(N938), .B0(N230), .Y(N952) );
  NAND2X2TF U233 ( .A(N580), .B(N357), .Y(N933) );
  AOI22XLTF U234 ( .A0(X_IN[2]), .A1(N818), .B0(X_IN[3]), .B1(N457), .Y(N437)
         );
  INVX2TF U235 ( .A(N986), .Y(N158) );
  AOI2BB1X2TF U236 ( .A0N(N980), .A1N(N979), .B0(N978), .Y(N1028) );
  OAI21XLTF U237 ( .A0(N616), .A1(N615), .B0(N614), .Y(N617) );
  INVXLTF U238 ( .A(N615), .Y(N582) );
  NOR3BX2TF U239 ( .AN(ALU_TYPE[2]), .B(ALU_TYPE[0]), .C(ALU_TYPE[1]), .Y(N272) );
  NOR3XLTF U240 ( .A(N130), .B(N927), .C(N989), .Y(N837) );
  NAND2X2TF U241 ( .A(N987), .B(N946), .Y(N927) );
  AOI21XLTF U242 ( .A0(N838), .A1(N386), .B0(N385), .Y(N388) );
  AOI21XLTF U243 ( .A0(N840), .A1(N839), .B0(N838), .Y(N846) );
  INVXLTF U244 ( .A(N838), .Y(N389) );
  NOR3BX4TF U245 ( .AN(N397), .B(N394), .C(N150), .Y(N526) );
  AOI21X2TF U246 ( .A0(N783), .A1(N319), .B0(N398), .Y(N394) );
  AOI222X4TF U247 ( .A0(XTEMP[9]), .A1(X_IN[9]), .B0(XTEMP[9]), .B1(N492), 
        .C0(X_IN[9]), .C1(N492), .Y(N501) );
  AOI222X4TF U248 ( .A0(N175), .A1(N502), .B0(N175), .B1(N478), .C0(N502), 
        .C1(N478), .Y(N492) );
  OAI31XLTF U249 ( .A0(OPER_A[1]), .A1(N933), .A2(OPER_A[0]), .B0(N848), .Y(
        N849) );
  OAI21X2TF U250 ( .A0(N527), .A1(N136), .B0(N257), .Y(OPER_A[1]) );
  NAND2X2TF U251 ( .A(N779), .B(N63), .Y(N574) );
  NOR2X4TF U252 ( .A(N398), .B(N785), .Y(N823) );
  AOI22XLTF U253 ( .A0(DIVISION_HEAD[5]), .A1(N115), .B0(X_IN[7]), .B1(N823), 
        .Y(N400) );
  AOI22XLTF U254 ( .A0(X_IN[10]), .A1(N155), .B0(X_IN[11]), .B1(N823), .Y(N439) );
  NOR4X2TF U255 ( .A(N733), .B(N960), .C(N378), .D(N377), .Y(N727) );
  NOR2X2TF U256 ( .A(N349), .B(N619), .Y(N581) );
  NOR2BX2TF U257 ( .AN(N559), .B(N395), .Y(N644) );
  INVX2TF U258 ( .A(N160), .Y(N161) );
  INVX2TF U259 ( .A(N160), .Y(N162) );
  AOI22X2TF U260 ( .A0(N356), .A1(N354), .B0(N957), .B1(N357), .Y(N939) );
  XNOR2X1TF U261 ( .A(OPER_A[12]), .B(ADD_X_132_1_N2), .Y(N163) );
  CMPR32X2TF U262 ( .A(OPER_A[7]), .B(OPER_B[7]), .C(ADD_X_132_1_N7), .CO(
        ADD_X_132_1_N6), .S(SUM_AB[7]) );
  CMPR32X2TF U263 ( .A(OPER_A[6]), .B(OPER_B[6]), .C(ADD_X_132_1_N8), .CO(
        ADD_X_132_1_N7), .S(SUM_AB[6]) );
  XNOR2X2TF U264 ( .A(N163), .B(OPER_B[12]), .Y(SUM_AB[12]) );
  INVX2TF U265 ( .A(OPER_A[0]), .Y(N842) );
  OAI21X2TF U266 ( .A0(N179), .A1(N136), .B0(N256), .Y(OPER_A[0]) );
  NOR2X1TF U267 ( .A(ALU_TYPE[2]), .B(ALU_TYPE[0]), .Y(N210) );
  AOI222XLTF U268 ( .A0(DIVISION_HEAD[1]), .A1(DIVISION_HEAD[0]), .B0(
        DIVISION_HEAD[1]), .B1(N325), .C0(DIVISION_HEAD[0]), .C1(N324), .Y(
        N327) );
  OAI31X1TF U269 ( .A0(N151), .A1(N966), .A2(N965), .B0(N964), .Y(N967) );
  AOI22X1TF U270 ( .A0(N130), .A1(N187), .B0(POST_WORK), .B1(N61), .Y(N255) );
  NAND2X1TF U271 ( .A(N324), .B(N742), .Y(N326) );
  NOR2X1TF U272 ( .A(SUM_AB[10]), .B(N500), .Y(N513) );
  NAND2X1TF U273 ( .A(N491), .B(N490), .Y(N500) );
  NOR2X1TF U274 ( .A(SUM_AB[8]), .B(N475), .Y(N491) );
  OA22X1TF U275 ( .A0(N785), .A1(N573), .B0(N780), .B1(N781), .Y(N319) );
  INVX2TF U276 ( .A(N946), .Y(N230) );
  OAI21X1TF U277 ( .A0(N965), .A1(N625), .B0(N732), .Y(N978) );
  NOR2X2TF U278 ( .A(N230), .B(N144), .Y(N921) );
  OR2X2TF U279 ( .A(N978), .B(N211), .Y(N946) );
  NOR2X1TF U280 ( .A(\INDEX[2] ), .B(N636), .Y(N322) );
  NAND2X1TF U281 ( .A(N129), .B(N128), .Y(N636) );
  OAI21X1TF U282 ( .A0(DIVISION_HEAD[12]), .A1(N564), .B0(N348), .Y(N965) );
  AOI2BB1X1TF U283 ( .A0N(DIVISION_HEAD[6]), .A1N(N337), .B0(Y_IN[6]), .Y(N335) );
  AOI21X1TF U284 ( .A0(N206), .A1(N527), .B0(N334), .Y(N337) );
  AOI2BB1X1TF U285 ( .A0N(DIVISION_HEAD[4]), .A1N(N333), .B0(Y_IN[4]), .Y(N331) );
  NAND2X1TF U286 ( .A(N929), .B(N921), .Y(N949) );
  AOI2BB1X1TF U287 ( .A0N(N623), .A1N(N353), .B0(N979), .Y(N211) );
  NOR2X1TF U288 ( .A(PRE_WORK), .B(N350), .Y(N352) );
  NAND2X1TF U289 ( .A(N122), .B(N177), .Y(N620) );
  NOR2X1TF U290 ( .A(N124), .B(N643), .Y(N350) );
  NAND2X1TF U291 ( .A(N106), .B(N272), .Y(N615) );
  NAND2X1TF U292 ( .A(N581), .B(N395), .Y(N625) );
  NOR2X1TF U293 ( .A(Y_IN[3]), .B(N734), .Y(N329) );
  NAND2X1TF U294 ( .A(N166), .B(N178), .Y(N349) );
  AOI211X1TF U295 ( .A0(N231), .A1(N623), .B0(N962), .C0(N622), .Y(N626) );
  NAND2X1TF U296 ( .A(N467), .B(N473), .Y(N485) );
  NAND2X2TF U297 ( .A(N562), .B(N397), .Y(N473) );
  CLKBUFX2TF U298 ( .A(N798), .Y(N205) );
  AOI211X1TF U299 ( .A0(Y_IN[11]), .A1(N315), .B0(Y_IN[12]), .C0(N296), .Y(
        N783) );
  NAND2X1TF U300 ( .A(N121), .B(N122), .Y(N973) );
  NAND3X1TF U301 ( .A(N979), .B(N151), .C(N615), .Y(N732) );
  AND2X2TF U302 ( .A(N106), .B(N159), .Y(N231) );
  NAND2X1TF U303 ( .A(N190), .B(N376), .Y(N358) );
  NAND2X1TF U304 ( .A(N124), .B(N322), .Y(N376) );
  NAND2X1TF U305 ( .A(N121), .B(N188), .Y(N619) );
  CLKBUFX2TF U306 ( .A(Y_IN[5]), .Y(N206) );
  AND2X2TF U307 ( .A(N210), .B(ALU_TYPE[1]), .Y(N232) );
  NOR3X1TF U308 ( .A(N621), .B(N620), .C(N793), .Y(N622) );
  OR3X1TF U309 ( .A(N899), .B(N898), .C(N225), .Y(N676) );
  OAI2BB2XLTF U310 ( .B0(N900), .B1(N989), .A0N(C152_DATA4_6), .A1N(N139), .Y(
        N225) );
  OAI2BB2XLTF U311 ( .B0(N897), .B1(N941), .A0N(N230), .A1N(OPER_B[6]), .Y(
        N898) );
  INVX2TF U312 ( .A(N473), .Y(N489) );
  AOI32X1TF U313 ( .A0(N987), .A1(N986), .A2(N985), .B0(N958), .B1(N986), .Y(
        N1036) );
  NAND2X1TF U314 ( .A(N581), .B(DP_OP_333_124_4748_N57), .Y(N406) );
  NAND2X1TF U315 ( .A(N977), .B(DP_OP_333_124_4748_N57), .Y(N736) );
  INVX2TF U316 ( .A(N375), .Y(N779) );
  NAND2X1TF U317 ( .A(N395), .B(N977), .Y(N375) );
  NOR2BX2TF U318 ( .AN(N562), .B(N572), .Y(N830) );
  NOR2X1TF U319 ( .A(N190), .B(N615), .Y(N363) );
  NAND2X1TF U320 ( .A(N921), .B(N888), .Y(N911) );
  NOR2X1TF U321 ( .A(N131), .B(N927), .Y(N923) );
  AOI21X1TF U322 ( .A0(N966), .A1(N984), .B0(N374), .Y(N987) );
  NAND2X1TF U323 ( .A(N166), .B(STEP[3]), .Y(N647) );
  NOR2X2TF U324 ( .A(N349), .B(N620), .Y(N977) );
  NAND2X1TF U325 ( .A(N350), .B(N190), .Y(N355) );
  NOR3BX1TF U326 ( .AN(ALU_TYPE[0]), .B(ALU_TYPE[1]), .C(ALU_TYPE[2]), .Y(N271) );
  AO22X1TF U327 ( .A0(N383), .A1(XTEMP[12]), .B0(N371), .B1(N982), .Y(N722) );
  AOI32X1TF U328 ( .A0(N984), .A1(N372), .A2(N975), .B0(N990), .B1(N372), .Y(
        N373) );
  NAND2X1TF U329 ( .A(N963), .B(DP_OP_333_124_4748_N57), .Y(N650) );
  NAND2X1TF U330 ( .A(N728), .B(N147), .Y(N630) );
  NAND2X1TF U331 ( .A(N139), .B(C152_DATA4_8), .Y(N226) );
  AOI32X1TF U332 ( .A0(N148), .A1(DIVISION_HEAD[4]), .A2(N766), .B0(N485), 
        .B1(DIVISION_HEAD[4]), .Y(N404) );
  OAI22X1TF U333 ( .A0(N544), .A1(N120), .B0(N502), .B1(N118), .Y(N503) );
  INVX2TF U334 ( .A(N1032), .Y(N1027) );
  OAI2BB2XLTF U335 ( .B0(N131), .B1(N989), .A0N(N989), .A1N(N131), .Y(N991) );
  NOR2X2TF U336 ( .A(N779), .B(N205), .Y(N777) );
  INVX2TF U337 ( .A(N146), .Y(N793) );
  OAI211X1TF U338 ( .A0(N977), .A1(N358), .B0(N582), .C0(N616), .Y(N359) );
  NAND2X1TF U339 ( .A(N732), .B(N117), .Y(N961) );
  NAND2X1TF U340 ( .A(N361), .B(N146), .Y(N559) );
  NOR2X1TF U341 ( .A(N973), .B(N647), .Y(N579) );
  NOR2X1TF U342 ( .A(N620), .B(N971), .Y(N580) );
  NAND2X1TF U343 ( .A(STEP[2]), .B(N178), .Y(N971) );
  INVX2TF U344 ( .A(N231), .Y(N979) );
  OAI32X1TF U345 ( .A0(N735), .A1(N192), .A2(N961), .B0(N734), .B1(N736), .Y(
        N694) );
  OAI21X1TF U346 ( .A0(N190), .A1(N733), .B0(N732), .Y(N695) );
  AOI22X1TF U347 ( .A0(N558), .A1(N130), .B0(N557), .B1(N556), .Y(N707) );
  INVX2TF U348 ( .A(N558), .Y(N556) );
  OAI31X1TF U349 ( .A0(N555), .A1(N554), .A2(N553), .B0(N552), .Y(N557) );
  AOI211X1TF U350 ( .A0(N551), .A1(XTEMP[12]), .B0(N550), .C0(N549), .Y(N552)
         );
  OAI31X1TF U351 ( .A0(DIVISION_HEAD[1]), .A1(N548), .A2(N176), .B0(N547), .Y(
        N551) );
  AOI22X1TF U352 ( .A0(N546), .A1(N545), .B0(XTEMP[11]), .B1(N829), .Y(N547)
         );
  OAI22X1TF U353 ( .A0(DIVISION_HEAD[0]), .A1(N544), .B0(DIVISION_REMA[8]), 
        .B1(N175), .Y(N545) );
  INVX2TF U354 ( .A(N554), .Y(N546) );
  NOR2X1TF U355 ( .A(XTEMP[11]), .B(N829), .Y(N548) );
  OAI22X1TF U356 ( .A0(DIVISION_HEAD[12]), .A1(N164), .B0(XTEMP[12]), .B1(N734), .Y(N553) );
  OAI21X1TF U357 ( .A0(XTEMP[11]), .A1(N829), .B0(N543), .Y(N554) );
  AOI22X1TF U358 ( .A0(DIVISION_HEAD[0]), .A1(N544), .B0(DIVISION_HEAD[1]), 
        .B1(N176), .Y(N543) );
  AOI21X1TF U359 ( .A0(DIVISION_HEAD[11]), .A1(N171), .B0(N542), .Y(N555) );
  AOI211X1TF U360 ( .A0(DIVISION_REMA[6]), .A1(N541), .B0(N540), .C0(N539), 
        .Y(N542) );
  NOR2X1TF U361 ( .A(DIVISION_HEAD[11]), .B(N171), .Y(N539) );
  AOI21X1TF U362 ( .A0(DIVISION_HEAD[9]), .A1(N170), .B0(N537), .Y(N538) );
  AOI211X1TF U363 ( .A0(DIVISION_REMA[4]), .A1(N536), .B0(N535), .C0(N534), 
        .Y(N537) );
  NOR2X1TF U364 ( .A(DIVISION_HEAD[9]), .B(N170), .Y(N534) );
  AOI21X1TF U365 ( .A0(DIVISION_HEAD[7]), .A1(N752), .B0(N532), .Y(N533) );
  AOI211X1TF U366 ( .A0(N531), .A1(DIVISION_REMA[2]), .B0(N530), .C0(N529), 
        .Y(N532) );
  NOR2X1TF U367 ( .A(DIVISION_HEAD[7]), .B(N752), .Y(N530) );
  OAI21X1TF U368 ( .A0(DIVISION_HEAD[5]), .A1(N184), .B0(N528), .Y(N531) );
  OAI211X1TF U369 ( .A0(DIVISION_REMA[1]), .A1(N527), .B0(DIVISION_REMA[0]), 
        .C0(N179), .Y(N528) );
  OAI21X1TF U370 ( .A0(N392), .A1(N187), .B0(N391), .Y(N720) );
  OAI22X1TF U371 ( .A0(N145), .A1(N389), .B0(N780), .B1(N655), .Y(N390) );
  OAI211X1TF U372 ( .A0(N384), .A1(N839), .B0(N627), .C0(N655), .Y(N385) );
  OAI21X1TF U373 ( .A0(N123), .A1(N969), .B0(N968), .Y(N670) );
  OAI21X1TF U374 ( .A0(N967), .A1(N987), .B0(N969), .Y(N968) );
  OR4X2TF U375 ( .A(N962), .B(N961), .C(N960), .D(N959), .Y(N969) );
  OAI22X1TF U376 ( .A0(N145), .A1(N957), .B0(N956), .B1(N990), .Y(N959) );
  OAI21X1TF U377 ( .A0(N612), .A1(N601), .B0(N600), .Y(N702) );
  AOI31X1TF U378 ( .A0(N599), .A1(N604), .A2(N606), .B0(N598), .Y(N601) );
  OAI22X1TF U379 ( .A0(N128), .A1(N597), .B0(N608), .B1(N604), .Y(N598) );
  AOI22X1TF U380 ( .A0(N612), .A1(N92), .B0(N596), .B1(N595), .Y(N703) );
  AOI211X1TF U381 ( .A0(N610), .A1(N182), .B0(N594), .C0(N807), .Y(N596) );
  AOI21X1TF U382 ( .A0(N593), .A1(N793), .B0(N194), .Y(N594) );
  OAI21X1TF U383 ( .A0(N128), .A1(N635), .B0(N634), .Y(N699) );
  AOI31X1TF U384 ( .A0(N633), .A1(N636), .A2(N632), .B0(N631), .Y(N634) );
  OAI32X1TF U385 ( .A0(N644), .A1(N645), .A2(N636), .B0(N632), .B1(N644), .Y(
        N631) );
  OAI21X1TF U386 ( .A0(N129), .A1(N635), .B0(N321), .Y(N726) );
  OAI21X1TF U387 ( .A0(N320), .A1(N394), .B0(N635), .Y(N321) );
  AOI32X1TF U388 ( .A0(N644), .A1(N650), .A2(N387), .B0(N182), .B1(N650), .Y(
        N320) );
  OAI31X1TF U389 ( .A0(N645), .A1(N644), .A2(N643), .B0(N642), .Y(N698) );
  AOI22X1TF U390 ( .A0(\INDEX[2] ), .A1(N641), .B0(N640), .B1(N639), .Y(N642)
         );
  OAI21X1TF U391 ( .A0(N638), .A1(N644), .B0(N637), .Y(N641) );
  OAI211X1TF U392 ( .A0(N145), .A1(N380), .B0(N730), .C0(N379), .Y(N721) );
  AOI22X1TF U393 ( .A0(STEP[3]), .A1(N727), .B0(N386), .B1(N589), .Y(N379) );
  NOR2X1TF U394 ( .A(N645), .B(N639), .Y(N637) );
  AOI21X1TF U395 ( .A0(\INDEX[2] ), .A1(N640), .B0(N387), .Y(N639) );
  INVX2TF U396 ( .A(N635), .Y(N645) );
  INVX2TF U397 ( .A(N632), .Y(N640) );
  OAI211X1TF U398 ( .A0(N193), .A1(N630), .B0(N646), .C0(N629), .Y(N700) );
  AOI21X1TF U399 ( .A0(N727), .A1(N177), .B0(N628), .Y(N629) );
  NOR3X1TF U400 ( .A(STEP[3]), .B(N145), .C(N619), .Y(N962) );
  AOI211X1TF U401 ( .A0(N840), .A1(N386), .B0(N383), .C0(N382), .Y(N627) );
  AOI21X1TF U402 ( .A0(N396), .A1(N381), .B0(N793), .Y(N382) );
  NOR2X1TF U403 ( .A(N144), .B(N839), .Y(N386) );
  OAI22X1TF U404 ( .A0(N90), .A1(N613), .B0(N612), .B1(N611), .Y(N701) );
  AOI21X1TF U405 ( .A0(\INDEX[2] ), .A1(N610), .B0(N609), .Y(N611) );
  OAI22X1TF U406 ( .A0(N608), .A1(N607), .B0(N606), .B1(N605), .Y(N609) );
  INVX2TF U407 ( .A(N603), .Y(N608) );
  AOI21X1TF U408 ( .A0(N604), .A1(N603), .B0(N602), .Y(N613) );
  OAI211X1TF U409 ( .A0(N731), .A1(N166), .B0(N730), .C0(N729), .Y(N696) );
  NOR2X1TF U410 ( .A(N735), .B(N373), .Y(N730) );
  OAI21X1TF U411 ( .A0(N361), .A1(N273), .B0(N103), .Y(N372) );
  INVX2TF U412 ( .A(N736), .Y(N735) );
  OAI22X1TF U413 ( .A0(N188), .A1(N971), .B0(N839), .B1(N984), .Y(N653) );
  AOI211X1TF U414 ( .A0(N727), .A1(N188), .B0(N652), .C0(N651), .Y(N656) );
  INVX2TF U415 ( .A(N274), .Y(N649) );
  AOI31X1TF U416 ( .A0(N973), .A1(N381), .A2(N396), .B0(N793), .Y(N274) );
  AOI21X1TF U417 ( .A0(N988), .A1(N618), .B0(N617), .Y(N646) );
  OAI22X1TF U418 ( .A0(N612), .A1(N592), .B0(N591), .B1(N203), .Y(N704) );
  AOI21X1TF U419 ( .A0(N607), .A1(N603), .B0(N602), .Y(N591) );
  OAI21X1TF U420 ( .A0(N90), .A1(N606), .B0(N599), .Y(N605) );
  INVX2TF U421 ( .A(N630), .Y(N599) );
  INVX2TF U422 ( .A(N612), .Y(N595) );
  OAI31X1TF U423 ( .A0(N621), .A1(N620), .A2(N793), .B0(N593), .Y(N603) );
  OAI32X1TF U424 ( .A0(N590), .A1(N840), .A2(N589), .B0(N958), .B1(N590), .Y(
        N593) );
  INVX2TF U425 ( .A(N588), .Y(N590) );
  AOI21X1TF U426 ( .A0(N610), .A1(N200), .B0(N587), .Y(N592) );
  AOI32X1TF U427 ( .A0(N581), .A1(N147), .A2(N193), .B0(N977), .B1(N146), .Y(
        N583) );
  AOI31X1TF U428 ( .A0(N103), .A1(N840), .A2(N839), .B0(N961), .Y(N584) );
  INVX2TF U429 ( .A(N597), .Y(N610) );
  AOI22X1TF U430 ( .A0(N920), .A1(N921), .B0(N230), .B1(OPER_B[8]), .Y(N227)
         );
  OAI21X1TF U431 ( .A0(N919), .A1(N185), .B0(N918), .Y(N920) );
  AOI211X1TF U432 ( .A0(N937), .A1(OPER_B[9]), .B0(N917), .C0(N916), .Y(N918)
         );
  OAI32X1TF U433 ( .A0(OPER_A[8]), .A1(N915), .A2(N933), .B0(N914), .B1(N913), 
        .Y(N916) );
  AOI21X1TF U434 ( .A0(N930), .A1(N915), .B0(N929), .Y(N913) );
  NOR3X1TF U435 ( .A(N928), .B(OPER_B[8]), .C(N912), .Y(N917) );
  AOI21X1TF U436 ( .A0(N912), .A1(N939), .B0(N938), .Y(N919) );
  OAI21X1TF U437 ( .A0(N463), .A1(N462), .B0(N473), .Y(N464) );
  AOI22X1TF U438 ( .A0(DIVISION_HEAD[11]), .A1(N116), .B0(X_IN[12]), .B1(N156), 
        .Y(N458) );
  AOI22X1TF U439 ( .A0(SUM_AB[6]), .A1(N153), .B0(N507), .B1(N1009), .Y(N460)
         );
  OAI22X1TF U440 ( .A0(N455), .A1(N120), .B0(N454), .B1(N118), .Y(N463) );
  OAI211X1TF U441 ( .A0(N1027), .A1(N1008), .B0(N1007), .C0(N1006), .Y(N664)
         );
  AOI22X1TF U442 ( .A0(DIVISION_HEAD[5]), .A1(N132), .B0(ZTEMP[5]), .B1(N158), 
        .Y(N1007) );
  OAI211X1TF U443 ( .A0(N1027), .A1(N1014), .B0(N1013), .C0(N1012), .Y(N662)
         );
  AOI22X1TF U444 ( .A0(DIVISION_HEAD[7]), .A1(N132), .B0(ZTEMP[7]), .B1(N158), 
        .Y(N1013) );
  OAI211X1TF U445 ( .A0(N1027), .A1(N1002), .B0(N1001), .C0(N1000), .Y(N666)
         );
  AOI22X1TF U446 ( .A0(DIVISION_HEAD[3]), .A1(N132), .B0(ZTEMP[3]), .B1(N1028), 
        .Y(N1001) );
  AOI22X1TF U447 ( .A0(SUM_AB[8]), .A1(N111), .B0(N1015), .B1(N1032), .Y(N1016) );
  AOI22X1TF U448 ( .A0(DIVISION_HEAD[8]), .A1(N133), .B0(ZTEMP[8]), .B1(N158), 
        .Y(N1017) );
  AOI22X1TF U449 ( .A0(SUM_AB[2]), .A1(N111), .B0(N997), .B1(N1032), .Y(N998)
         );
  AOI22X1TF U450 ( .A0(DIVISION_HEAD[2]), .A1(N133), .B0(ZTEMP[2]), .B1(N158), 
        .Y(N999) );
  AOI22X1TF U451 ( .A0(SUM_AB[4]), .A1(N111), .B0(N1003), .B1(N1032), .Y(N1004) );
  AOI22X1TF U452 ( .A0(DIVISION_HEAD[4]), .A1(N133), .B0(ZTEMP[4]), .B1(N158), 
        .Y(N1005) );
  AOI22X1TF U453 ( .A0(SUM_AB[1]), .A1(N111), .B0(N994), .B1(N1032), .Y(N995)
         );
  AOI22X1TF U454 ( .A0(DIVISION_HEAD[1]), .A1(N133), .B0(ZTEMP[1]), .B1(N158), 
        .Y(N996) );
  AOI22X1TF U455 ( .A0(SUM_AB[6]), .A1(N111), .B0(N1009), .B1(N1032), .Y(N1010) );
  AOI22X1TF U456 ( .A0(DIVISION_HEAD[6]), .A1(N133), .B0(ZTEMP[6]), .B1(N158), 
        .Y(N1011) );
  OAI211X1TF U457 ( .A0(N1027), .A1(N1020), .B0(N1019), .C0(N1018), .Y(N660)
         );
  AOI22X1TF U458 ( .A0(DIVISION_HEAD[9]), .A1(N132), .B0(ZTEMP[9]), .B1(N1028), 
        .Y(N1019) );
  INVX2TF U459 ( .A(N899), .Y(N222) );
  AOI31X1TF U460 ( .A0(N853), .A1(N852), .A2(N851), .B0(N941), .Y(N855) );
  AOI32X1TF U461 ( .A0(N850), .A1(OPER_B[2]), .A2(N939), .B0(N938), .B1(
        OPER_B[2]), .Y(N851) );
  AOI22X1TF U462 ( .A0(N937), .A1(OPER_B[3]), .B0(OPER_A[2]), .B1(N849), .Y(
        N852) );
  AOI31X1TF U463 ( .A0(N939), .A1(N181), .A2(N845), .B0(N844), .Y(N853) );
  AOI211X1TF U464 ( .A0(N843), .A1(N842), .B0(OPER_A[2]), .C0(N933), .Y(N844)
         );
  AOI211X1TF U465 ( .A0(N230), .A1(OPER_B[10]), .B0(N944), .C0(N945), .Y(N228)
         );
  AOI21X1TF U466 ( .A0(N992), .A1(N989), .B0(N927), .Y(N945) );
  AOI21X1TF U467 ( .A0(N943), .A1(N942), .B0(N941), .Y(N944) );
  AOI32X1TF U468 ( .A0(N940), .A1(OPER_B[10]), .A2(N939), .B0(N938), .B1(
        OPER_B[10]), .Y(N942) );
  AOI211X1TF U469 ( .A0(N937), .A1(OPER_B[11]), .B0(N936), .C0(N935), .Y(N943)
         );
  OAI32X1TF U470 ( .A0(OPER_A[10]), .A1(N934), .A2(N933), .B0(N932), .B1(N931), 
        .Y(N935) );
  AOI21X1TF U471 ( .A0(N930), .A1(N934), .B0(N929), .Y(N931) );
  NOR3X1TF U472 ( .A(N928), .B(OPER_B[10]), .C(N940), .Y(N936) );
  OAI22X1TF U473 ( .A0(N489), .A1(N488), .B0(N487), .B1(N175), .Y(N711) );
  AOI211X1TF U474 ( .A0(N1015), .A1(N507), .B0(N484), .C0(N483), .Y(N488) );
  OAI211X1TF U475 ( .A0(N482), .A1(N624), .B0(N481), .C0(N480), .Y(N483) );
  AOI22X1TF U476 ( .A0(XTEMP[9]), .A1(N116), .B0(N816), .B1(SUM_AB[12]), .Y(
        N480) );
  NOR2X1TF U477 ( .A(DIVISION_HEAD[12]), .B(N486), .Y(N479) );
  AOI22X1TF U478 ( .A0(X_IN[8]), .A1(N478), .B0(INTADD_0_N1), .B1(N502), .Y(
        N486) );
  OAI22X1TF U479 ( .A0(N477), .A1(N120), .B0(N476), .B1(N118), .Y(N484) );
  AOI211X1TF U480 ( .A0(OPER_B[6]), .A1(N896), .B0(N895), .C0(N894), .Y(N897)
         );
  OAI32X1TF U481 ( .A0(OPER_A[6]), .A1(N893), .A2(N933), .B0(N892), .B1(N891), 
        .Y(N894) );
  AOI21X1TF U482 ( .A0(N930), .A1(N893), .B0(N929), .Y(N891) );
  INVX2TF U483 ( .A(N933), .Y(N930) );
  OAI31X1TF U484 ( .A0(N928), .A1(OPER_B[6]), .A2(N890), .B0(N889), .Y(N895)
         );
  AOI21X1TF U485 ( .A0(OPER_B[7]), .A1(N888), .B0(N887), .Y(N889) );
  OAI21X1TF U486 ( .A0(N928), .A1(N886), .B0(N885), .Y(N896) );
  AOI32X1TF U487 ( .A0(N405), .A1(N404), .A2(N403), .B0(N489), .B1(N404), .Y(
        N719) );
  OAI211X1TF U488 ( .A0(N401), .A1(N574), .B0(N400), .C0(N399), .Y(N402) );
  AOI22X1TF U489 ( .A0(X_IN[6]), .A1(N156), .B0(X_IN[5]), .B1(N126), .Y(N399)
         );
  AOI22X1TF U490 ( .A0(DIVISION_HEAD[3]), .A1(N751), .B0(SUM_AB[0]), .B1(N393), 
        .Y(N405) );
  AOI32X1TF U491 ( .A0(N424), .A1(N473), .A2(N423), .B0(N489), .B1(N167), .Y(
        N717) );
  AOI211X1TF U492 ( .A0(DIVISION_HEAD[7]), .A1(N116), .B0(N422), .C0(N421), 
        .Y(N423) );
  OAI211X1TF U493 ( .A0(N118), .A1(N766), .B0(N420), .C0(N419), .Y(N421) );
  AOI21X1TF U494 ( .A0(N507), .A1(N997), .B0(N418), .Y(N419) );
  OAI22X1TF U495 ( .A0(N527), .A1(N119), .B0(N167), .B1(N467), .Y(N418) );
  AOI22X1TF U496 ( .A0(X_IN[1]), .A1(N457), .B0(N816), .B1(SUM_AB[6]), .Y(N420) );
  OAI21X1TF U497 ( .A0(N514), .A1(N765), .B0(N415), .Y(N422) );
  AOI22X1TF U498 ( .A0(X_IN[8]), .A1(N156), .B0(X_IN[7]), .B1(N126), .Y(N415)
         );
  AOI32X1TF U499 ( .A0(N443), .A1(N473), .A2(N442), .B0(N489), .B1(N536), .Y(
        N715) );
  AOI211X1TF U500 ( .A0(N507), .A1(N1003), .B0(N441), .C0(N440), .Y(N442) );
  AOI22X1TF U501 ( .A0(DIVISION_HEAD[9]), .A1(N115), .B0(X_IN[9]), .B1(N126), 
        .Y(N438) );
  OAI22X1TF U502 ( .A0(N168), .A1(N120), .B0(N536), .B1(N467), .Y(N441) );
  AOI32X1TF U503 ( .A0(N474), .A1(N473), .A2(N472), .B0(N489), .B1(N477), .Y(
        N712) );
  OAI211X1TF U504 ( .A0(N520), .A1(N1014), .B0(N469), .C0(N468), .Y(N470) );
  AOI22X1TF U505 ( .A0(DIVISION_HEAD[12]), .A1(N115), .B0(X_IN[12]), .B1(N125), 
        .Y(N468) );
  AOI22X1TF U506 ( .A0(DIVISION_HEAD[11]), .A1(N822), .B0(DIVISION_HEAD[10]), 
        .B1(N150), .Y(N469) );
  OAI22X1TF U507 ( .A0(N476), .A1(N624), .B0(N574), .B1(N512), .Y(N471) );
  AOI32X1TF U508 ( .A0(N414), .A1(N473), .A2(N413), .B0(N489), .B1(N527), .Y(
        N718) );
  AOI211X1TF U509 ( .A0(N507), .A1(N994), .B0(N412), .C0(N411), .Y(N413) );
  OAI211X1TF U510 ( .A0(N574), .A1(N444), .B0(N410), .C0(N409), .Y(N411) );
  AOI21X1TF U511 ( .A0(DIVISION_HEAD[4]), .A1(N751), .B0(N408), .Y(N409) );
  OAI22X1TF U512 ( .A0(N527), .A1(N467), .B0(N766), .B1(N624), .Y(N408) );
  AOI22X1TF U513 ( .A0(DIVISION_HEAD[6]), .A1(N116), .B0(X_IN[7]), .B1(N155), 
        .Y(N410) );
  OAI22X1TF U514 ( .A0(N476), .A1(N407), .B0(N502), .B1(N765), .Y(N412) );
  OAI22X1TF U515 ( .A0(N526), .A1(N499), .B0(N498), .B1(N544), .Y(N710) );
  AOI211X1TF U516 ( .A0(SUM_AB[9]), .A1(N154), .B0(N496), .C0(N495), .Y(N499)
         );
  OAI211X1TF U517 ( .A0(N1020), .A1(N520), .B0(N494), .C0(N493), .Y(N495) );
  AOI22X1TF U518 ( .A0(XTEMP[10]), .A1(N116), .B0(X_IN[7]), .B1(N818), .Y(N494) );
  OAI22X1TF U519 ( .A0(N175), .A1(N120), .B0(N502), .B1(N624), .Y(N496) );
  AOI22X1TF U520 ( .A0(N205), .A1(N164), .B0(N797), .B1(N796), .Y(N686) );
  AOI211X1TF U521 ( .A0(DIVISION_REMA[7]), .A1(N751), .B0(N795), .C0(N794), 
        .Y(N797) );
  OAI211X1TF U522 ( .A0(N172), .A1(N793), .B0(N792), .C0(N791), .Y(N794) );
  AOI22X1TF U523 ( .A0(N790), .A1(N789), .B0(N1015), .B1(N813), .Y(N791) );
  AOI21X1TF U524 ( .A0(SUM_AB[8]), .A1(N475), .B0(N491), .Y(N1015) );
  AOI32X1TF U525 ( .A0(N788), .A1(N787), .A2(N786), .B0(N785), .B1(N787), .Y(
        N789) );
  OAI32X1TF U526 ( .A0(N784), .A1(N783), .A2(X_IN[0]), .B0(N782), .B1(N784), 
        .Y(N787) );
  AOI22X1TF U527 ( .A0(DIVISION_REMA[8]), .A1(N779), .B0(SUM_AB[8]), .B1(N161), 
        .Y(N792) );
  AOI22X1TF U528 ( .A0(SUM_AB[10]), .A1(N112), .B0(N1021), .B1(N1032), .Y(
        N1022) );
  AOI22X1TF U529 ( .A0(DIVISION_HEAD[10]), .A1(N133), .B0(ZTEMP[10]), .B1(N158), .Y(N1023) );
  AOI22X1TF U530 ( .A0(N489), .A1(N455), .B0(N453), .B1(N473), .Y(N714) );
  AOI21X1TF U531 ( .A0(DIVISION_HEAD[8]), .A1(N150), .B0(N446), .Y(N447) );
  OAI22X1TF U532 ( .A0(N455), .A1(N467), .B0(N520), .B1(N1008), .Y(N446) );
  AOI22X1TF U533 ( .A0(DIVISION_HEAD[10]), .A1(N115), .B0(X_IN[10]), .B1(N125), 
        .Y(N449) );
  OAI22X1TF U534 ( .A0(N454), .A1(N624), .B0(N574), .B1(N490), .Y(N452) );
  AOI32X1TF U535 ( .A0(N815), .A1(N832), .A2(N814), .B0(N830), .B1(N165), .Y(
        N684) );
  AOI21X1TF U536 ( .A0(N813), .A1(N1021), .B0(N812), .Y(N814) );
  AOI22X1TF U537 ( .A0(X_IN[2]), .A1(N126), .B0(X_IN[4]), .B1(N823), .Y(N808)
         );
  AOI22X1TF U538 ( .A0(DIVISION_HEAD[0]), .A1(N150), .B0(DIVISION_HEAD[1]), 
        .B1(N822), .Y(N809) );
  AOI22X1TF U539 ( .A0(Y_IN[10]), .A1(N807), .B0(X_IN[3]), .B1(N156), .Y(N810)
         );
  AOI22X1TF U540 ( .A0(N816), .A1(SUM_AB[1]), .B0(SUM_AB[10]), .B1(N162), .Y(
        N815) );
  OAI22X1TF U541 ( .A0(N526), .A1(N510), .B0(N509), .B1(N176), .Y(N709) );
  AOI21X1TF U542 ( .A0(N507), .A1(N1021), .B0(N506), .Y(N510) );
  OAI211X1TF U543 ( .A0(N514), .A1(N624), .B0(N505), .C0(N504), .Y(N506) );
  AOI22X1TF U544 ( .A0(XTEMP[11]), .A1(N116), .B0(SUM_AB[10]), .B1(N153), .Y(
        N505) );
  AOI21X1TF U545 ( .A0(SUM_AB[10]), .A1(N500), .B0(N513), .Y(N1021) );
  AOI32X1TF U546 ( .A0(N434), .A1(N473), .A2(N433), .B0(N489), .B1(N168), .Y(
        N716) );
  AOI211X1TF U547 ( .A0(DIVISION_HEAD[8]), .A1(N116), .B0(N432), .C0(N431), 
        .Y(N433) );
  OAI211X1TF U548 ( .A0(N574), .A1(N465), .B0(N430), .C0(N429), .Y(N431) );
  AOI21X1TF U549 ( .A0(DIVISION_HEAD[6]), .A1(N751), .B0(N428), .Y(N429) );
  OAI22X1TF U550 ( .A0(N168), .A1(N467), .B0(N520), .B1(N1002), .Y(N428) );
  OAI21X1TF U551 ( .A0(N515), .A1(N765), .B0(N425), .Y(N432) );
  AOI22X1TF U552 ( .A0(X_IN[8]), .A1(N126), .B0(X_IN[9]), .B1(N156), .Y(N425)
         );
  OAI211X1TF U553 ( .A0(N1027), .A1(N1026), .B0(N1025), .C0(N1024), .Y(N658)
         );
  AOI22X1TF U554 ( .A0(DIVISION_HEAD[11]), .A1(N133), .B0(ZTEMP[11]), .B1(N158), .Y(N1025) );
  OAI21X1TF U555 ( .A0(N777), .A1(N193), .B0(N578), .Y(N705) );
  OAI22X1TF U556 ( .A0(N577), .A1(N576), .B0(N779), .B1(N796), .Y(N578) );
  AOI22X1TF U557 ( .A0(Y_IN[0]), .A1(N807), .B0(DIVISION_REMA[1]), .B1(N146), 
        .Y(N575) );
  AOI21X1TF U558 ( .A0(N145), .A1(N736), .B0(N993), .Y(N577) );
  INVX2TF U559 ( .A(SUM_AB[0]), .Y(N993) );
  OAI22X1TF U560 ( .A0(N205), .A1(N740), .B0(N777), .B1(N184), .Y(N693) );
  AOI21X1TF U561 ( .A0(SUM_AB[1]), .A1(N162), .B0(N739), .Y(N740) );
  AOI22X1TF U562 ( .A0(DIVISION_REMA[0]), .A1(N751), .B0(N813), .B1(N994), .Y(
        N737) );
  AOI21X1TF U563 ( .A0(SUM_AB[1]), .A1(SUM_AB[0]), .B0(N416), .Y(N994) );
  AOI22X1TF U564 ( .A0(Y_IN[1]), .A1(N807), .B0(DIVISION_REMA[2]), .B1(N147), 
        .Y(N738) );
  OAI211X1TF U565 ( .A0(N1036), .A1(N1035), .B0(N1034), .C0(N1033), .Y(N657)
         );
  AOI32X1TF U566 ( .A0(N1035), .A1(N1032), .A2(N1031), .B0(N1030), .B1(N1032), 
        .Y(N1033) );
  AOI211X4TF U567 ( .A0(N992), .A1(N991), .B0(N990), .C0(N1028), .Y(N1032) );
  INVX2TF U568 ( .A(N987), .Y(N990) );
  AOI22X1TF U569 ( .A0(DIVISION_HEAD[12]), .A1(N133), .B0(ZTEMP[12]), .B1(
        N1028), .Y(N1034) );
  OAI31X1TF U570 ( .A0(N984), .A1(N131), .A2(N989), .B0(N983), .Y(N985) );
  AOI31X1TF U571 ( .A0(N192), .A1(N131), .A2(N982), .B0(N981), .Y(N983) );
  INVX2TF U572 ( .A(N1028), .Y(N986) );
  AOI31X1TF U573 ( .A0(N977), .A1(N976), .A2(N975), .B0(N974), .Y(N980) );
  OAI31X1TF U574 ( .A0(N973), .A1(N972), .A2(N971), .B0(N970), .Y(N974) );
  OAI22X1TF U575 ( .A0(N205), .A1(N769), .B0(N777), .B1(N174), .Y(N688) );
  AOI211X1TF U576 ( .A0(N1009), .A1(N813), .B0(N768), .C0(N767), .Y(N769) );
  OAI211X1TF U577 ( .A0(N766), .A1(N765), .B0(N773), .C0(N764), .Y(N767) );
  AOI22X1TF U578 ( .A0(DIVISION_REMA[7]), .A1(N146), .B0(SUM_AB[6]), .B1(N161), 
        .Y(N764) );
  INVX2TF U579 ( .A(N823), .Y(N765) );
  OAI21X1TF U580 ( .A0(N214), .A1(N118), .B0(N762), .Y(N768) );
  AOI22X1TF U581 ( .A0(Y_IN[6]), .A1(N807), .B0(DIVISION_REMA[5]), .B1(N751), 
        .Y(N762) );
  AOI21X1TF U582 ( .A0(SUM_AB[6]), .A1(N456), .B0(N466), .Y(N1009) );
  OAI22X1TF U583 ( .A0(N205), .A1(N757), .B0(N777), .B1(N173), .Y(N690) );
  AOI211X1TF U584 ( .A0(SUM_AB[4]), .A1(N162), .B0(N756), .C0(N755), .Y(N757)
         );
  OAI211X1TF U585 ( .A0(N754), .A1(N118), .B0(N773), .C0(N753), .Y(N755) );
  AOI22X1TF U586 ( .A0(DIVISION_REMA[5]), .A1(N147), .B0(N813), .B1(N1003), 
        .Y(N753) );
  AOI21X1TF U587 ( .A0(SUM_AB[4]), .A1(N435), .B0(N445), .Y(N1003) );
  OAI22X1TF U588 ( .A0(N214), .A1(N820), .B0(N752), .B1(N120), .Y(N756) );
  OAI22X1TF U589 ( .A0(N205), .A1(N745), .B0(N777), .B1(N180), .Y(N692) );
  AOI211X1TF U590 ( .A0(SUM_AB[2]), .A1(N162), .B0(N744), .C0(N743), .Y(N745)
         );
  OAI211X1TF U591 ( .A0(N742), .A1(N118), .B0(N773), .C0(N741), .Y(N743) );
  AOI22X1TF U592 ( .A0(DIVISION_REMA[3]), .A1(N147), .B0(N813), .B1(N997), .Y(
        N741) );
  AOI21X1TF U593 ( .A0(SUM_AB[2]), .A1(N417), .B0(N427), .Y(N997) );
  NOR2X1TF U594 ( .A(SUM_AB[0]), .B(SUM_AB[1]), .Y(N416) );
  OAI22X1TF U595 ( .A0(N754), .A1(N820), .B0(N184), .B1(N120), .Y(N744) );
  INVX2TF U596 ( .A(N939), .Y(N928) );
  OAI22X1TF U597 ( .A0(N526), .A1(N525), .B0(N524), .B1(N169), .Y(N708) );
  OAI21X1TF U598 ( .A0(N520), .A1(N1026), .B0(N519), .Y(N521) );
  AOI211X1TF U599 ( .A0(SUM_AB[11]), .A1(N153), .B0(N517), .C0(N516), .Y(N519)
         );
  OAI22X1TF U600 ( .A0(N176), .A1(N119), .B0(N514), .B1(N117), .Y(N517) );
  INVX2TF U601 ( .A(N507), .Y(N520) );
  OAI21X1TF U602 ( .A0(N777), .A1(N171), .B0(N776), .Y(N687) );
  OAI21X1TF U603 ( .A0(N775), .A1(N774), .B0(N796), .Y(N776) );
  INVX2TF U604 ( .A(N205), .Y(N796) );
  OAI211X1TF U605 ( .A0(N164), .A1(N793), .B0(N773), .C0(N772), .Y(N774) );
  AOI22X1TF U606 ( .A0(DIVISION_REMA[6]), .A1(N751), .B0(SUM_AB[7]), .B1(N161), 
        .Y(N772) );
  OAI211X1TF U607 ( .A0(N826), .A1(N1014), .B0(N771), .C0(N770), .Y(N775) );
  AOI22X1TF U608 ( .A0(X_IN[1]), .A1(N823), .B0(X_IN[0]), .B1(N156), .Y(N770)
         );
  OAI21X1TF U609 ( .A0(N466), .A1(N465), .B0(N475), .Y(N1014) );
  OAI22X1TF U610 ( .A0(N205), .A1(N761), .B0(N777), .B1(N170), .Y(N689) );
  AOI211X1TF U611 ( .A0(SUM_AB[5]), .A1(N162), .B0(N760), .C0(N759), .Y(N761)
         );
  OAI211X1TF U612 ( .A0(N826), .A1(N1008), .B0(N773), .C0(N758), .Y(N759) );
  OAI21X1TF U613 ( .A0(N445), .A1(N444), .B0(N456), .Y(N1008) );
  INVX2TF U614 ( .A(N820), .Y(N807) );
  OAI22X1TF U615 ( .A0(N205), .A1(N750), .B0(N777), .B1(N752), .Y(N691) );
  AOI211X1TF U616 ( .A0(SUM_AB[3]), .A1(N162), .B0(N749), .C0(N748), .Y(N750)
         );
  OAI211X1TF U617 ( .A0(N826), .A1(N1002), .B0(N773), .C0(N747), .Y(N748) );
  AOI222X4TF U618 ( .A0(N783), .A1(N125), .B0(N781), .B1(N155), .C0(N573), 
        .C1(N823), .Y(N773) );
  OAI21X1TF U619 ( .A0(N427), .A1(N426), .B0(N435), .Y(N1002) );
  OAI22X1TF U620 ( .A0(N746), .A1(N820), .B0(N180), .B1(N120), .Y(N749) );
  NOR3X1TF U621 ( .A(N790), .B(N150), .C(N572), .Y(N798) );
  AOI32X1TF U622 ( .A0(N806), .A1(N832), .A2(N805), .B0(N830), .B1(N172), .Y(
        N685) );
  OAI211X1TF U623 ( .A0(N826), .A1(N1020), .B0(N802), .C0(N801), .Y(N803) );
  AOI22X1TF U624 ( .A0(DIVISION_HEAD[1]), .A1(N147), .B0(X_IN[1]), .B1(N125), 
        .Y(N801) );
  OAI21X1TF U625 ( .A0(N491), .A1(N490), .B0(N500), .Y(N1020) );
  OAI21X1TF U626 ( .A0(N800), .A1(N820), .B0(N799), .Y(N804) );
  AOI22X1TF U627 ( .A0(DIVISION_REMA[8]), .A1(N150), .B0(N816), .B1(SUM_AB[0]), 
        .Y(N799) );
  AOI22X1TF U628 ( .A0(DIVISION_HEAD[0]), .A1(N822), .B0(SUM_AB[9]), .B1(N162), 
        .Y(N806) );
  OAI22X1TF U629 ( .A0(N526), .A1(N370), .B0(N369), .B1(N368), .Y(N723) );
  AOI211X1TF U630 ( .A0(N507), .A1(N1030), .B0(N366), .C0(N365), .Y(N370) );
  OAI31X1TF U631 ( .A0(XTEMP[12]), .A1(N367), .A2(N522), .B0(N364), .Y(N365)
         );
  INVX2TF U632 ( .A(N624), .Y(N457) );
  NAND2X2TF U633 ( .A(MODE_TYPE[1]), .B(N363), .Y(N624) );
  INVX2TF U634 ( .A(INTADD_0_N1), .Y(N478) );
  NOR2X1TF U635 ( .A(N179), .B(N766), .Y(INTADD_0_CI) );
  INVX2TF U636 ( .A(X_IN[0]), .Y(N766) );
  OAI22X1TF U637 ( .A0(N145), .A1(N1035), .B0(N515), .B1(N118), .Y(N366) );
  NOR2X2TF U638 ( .A(N406), .B(N1035), .Y(N507) );
  AOI31X1TF U639 ( .A0(N103), .A1(N130), .A2(N579), .B0(N360), .Y(N397) );
  OAI211X1TF U640 ( .A0(N130), .A1(N387), .B0(N371), .C0(N359), .Y(N360) );
  NOR2X1TF U641 ( .A(PRE_WORK), .B(N376), .Y(N618) );
  NOR2X1TF U642 ( .A(N383), .B(N961), .Y(N371) );
  INVX2TF U643 ( .A(N406), .Y(N383) );
  INVX2TF U644 ( .A(N633), .Y(N387) );
  AOI32X1TF U645 ( .A0(N833), .A1(N832), .A2(N831), .B0(N830), .B1(N829), .Y(
        N683) );
  AOI211X1TF U646 ( .A0(DIVISION_HEAD[3]), .A1(N147), .B0(N828), .C0(N827), 
        .Y(N831) );
  OAI211X1TF U647 ( .A0(N826), .A1(N1026), .B0(N825), .C0(N824), .Y(N827) );
  AOI22X1TF U648 ( .A0(X_IN[3]), .A1(N125), .B0(X_IN[5]), .B1(N823), .Y(N824)
         );
  AOI22X1TF U649 ( .A0(DIVISION_HEAD[1]), .A1(N150), .B0(DIVISION_HEAD[2]), 
        .B1(N822), .Y(N825) );
  OAI21X1TF U650 ( .A0(N513), .A1(N512), .B0(N1031), .Y(N1026) );
  INVX2TF U651 ( .A(N813), .Y(N826) );
  OAI21X1TF U652 ( .A0(N821), .A1(N820), .B0(N819), .Y(N828) );
  INVX2TF U653 ( .A(N117), .Y(N818) );
  INVX2TF U654 ( .A(N830), .Y(N832) );
  AOI22X1TF U655 ( .A0(N816), .A1(SUM_AB[2]), .B0(SUM_AB[11]), .B1(N162), .Y(
        N833) );
  OAI21X1TF U656 ( .A0(N830), .A1(N571), .B0(N570), .Y(N706) );
  OAI21X1TF U657 ( .A0(N830), .A1(N822), .B0(DIVISION_HEAD[3]), .Y(N570) );
  INVX2TF U658 ( .A(N467), .Y(N822) );
  AOI211X1TF U659 ( .A0(DIVISION_HEAD[2]), .A1(N150), .B0(N569), .C0(N568), 
        .Y(N571) );
  AOI22X1TF U660 ( .A0(N816), .A1(SUM_AB[3]), .B0(N1030), .B1(N813), .Y(N565)
         );
  NOR2X2TF U661 ( .A(N1035), .B(N736), .Y(N813) );
  NOR2X1TF U662 ( .A(N1035), .B(N1031), .Y(N1030) );
  INVX2TF U663 ( .A(SUM_AB[11]), .Y(N512) );
  INVX2TF U664 ( .A(SUM_AB[9]), .Y(N490) );
  INVX2TF U665 ( .A(SUM_AB[7]), .Y(N465) );
  NOR2X1TF U666 ( .A(SUM_AB[6]), .B(N456), .Y(N466) );
  INVX2TF U667 ( .A(SUM_AB[5]), .Y(N444) );
  NOR2X1TF U668 ( .A(SUM_AB[4]), .B(N435), .Y(N445) );
  INVX2TF U669 ( .A(SUM_AB[3]), .Y(N426) );
  NOR3X1TF U670 ( .A(SUM_AB[0]), .B(SUM_AB[2]), .C(SUM_AB[1]), .Y(N427) );
  INVX2TF U671 ( .A(SUM_AB[12]), .Y(N1035) );
  INVX2TF U672 ( .A(N574), .Y(N816) );
  AOI22X1TF U673 ( .A0(N103), .A1(SUM_AB[12]), .B0(X_IN[5]), .B1(N156), .Y(
        N566) );
  OAI21X1TF U674 ( .A0(N368), .A1(N137), .B0(N269), .Y(OPER_A[12]) );
  AOI22X1TF U675 ( .A0(X_IN[4]), .A1(N126), .B0(X_IN[6]), .B1(N823), .Y(N567)
         );
  AND2X2TF U676 ( .A(N780), .B(N785), .Y(N782) );
  INVX2TF U677 ( .A(N398), .Y(N790) );
  OAI22X1TF U678 ( .A0(N564), .A1(N820), .B0(N563), .B1(N118), .Y(N569) );
  NAND2X2TF U679 ( .A(N363), .B(N323), .Y(N820) );
  AOI32X1TF U680 ( .A0(N103), .A1(N131), .A2(N579), .B0(N633), .B1(N130), .Y(
        N560) );
  INVX2TF U681 ( .A(N363), .Y(N655) );
  AOI31X1TF U682 ( .A0(N122), .A1(N396), .A2(N395), .B0(N394), .Y(N562) );
  INVX2TF U683 ( .A(N318), .Y(N781) );
  OAI211X1TF U684 ( .A0(X_IN[12]), .A1(N563), .B0(N317), .C0(N316), .Y(N318)
         );
  OAI22X1TF U685 ( .A0(Y_IN[10]), .A1(N315), .B0(N314), .B1(N313), .Y(N316) );
  OAI22X1TF U686 ( .A0(X_IN[10]), .A1(N312), .B0(X_IN[11]), .B1(N800), .Y(N313) );
  OAI21X1TF U687 ( .A0(Y_IN[9]), .A1(N311), .B0(Y_IN[8]), .Y(N312) );
  AOI211X1TF U688 ( .A0(X_IN[10]), .A1(N778), .B0(N310), .C0(N309), .Y(N314)
         );
  AOI21X1TF U689 ( .A0(Y_IN[7]), .A1(N514), .B0(N308), .Y(N309) );
  AOI211X1TF U690 ( .A0(X_IN[8]), .A1(N307), .B0(N306), .C0(N305), .Y(N308) );
  NOR2X1TF U691 ( .A(Y_IN[7]), .B(N514), .Y(N306) );
  AOI21X1TF U692 ( .A0(N206), .A1(N482), .B0(N304), .Y(N307) );
  AOI211X1TF U693 ( .A0(X_IN[6]), .A1(N303), .B0(N302), .C0(N301), .Y(N304) );
  NOR2X1TF U694 ( .A(N206), .B(N482), .Y(N302) );
  AOI32X1TF U695 ( .A0(N300), .A1(N299), .A2(N326), .B0(N298), .B1(N299), .Y(
        N303) );
  OAI22X1TF U696 ( .A0(X_IN[4]), .A1(N754), .B0(N127), .B1(N746), .Y(N298) );
  OAI32X1TF U697 ( .A0(N297), .A1(N114), .A2(N324), .B0(X_IN[2]), .B1(N297), 
        .Y(N300) );
  INVX2TF U698 ( .A(X_IN[7]), .Y(N482) );
  INVX2TF U699 ( .A(X_IN[9]), .Y(N514) );
  NOR2X1TF U700 ( .A(Y_IN[9]), .B(N311), .Y(N310) );
  INVX2TF U701 ( .A(X_IN[11]), .Y(N311) );
  NOR2X1TF U702 ( .A(Y_IN[12]), .B(Y_IN[11]), .Y(N317) );
  INVX2TF U703 ( .A(N786), .Y(N573) );
  OR2X2TF U704 ( .A(MODE_TYPE[0]), .B(N323), .Y(N785) );
  INVX2TF U705 ( .A(MODE_TYPE[1]), .Y(N323) );
  OAI31X1TF U706 ( .A0(N293), .A1(N292), .A2(N291), .B0(N290), .Y(N294) );
  NOR2X1TF U707 ( .A(X_IN[10]), .B(N800), .Y(N291) );
  AOI211X1TF U708 ( .A0(X_IN[10]), .A1(N800), .B0(X_IN[9]), .C0(N778), .Y(N292) );
  AOI211X1TF U709 ( .A0(X_IN[9]), .A1(N778), .B0(N289), .C0(N288), .Y(N293) );
  AOI21X1TF U710 ( .A0(Y_IN[7]), .A1(N502), .B0(N287), .Y(N288) );
  AOI211X1TF U711 ( .A0(N286), .A1(X_IN[7]), .B0(N285), .C0(N284), .Y(N287) );
  NOR2X1TF U712 ( .A(Y_IN[7]), .B(N502), .Y(N285) );
  AOI21X1TF U713 ( .A0(N206), .A1(N476), .B0(N283), .Y(N286) );
  AOI211X1TF U714 ( .A0(N282), .A1(X_IN[5]), .B0(N281), .C0(N280), .Y(N283) );
  NOR2X1TF U715 ( .A(N206), .B(N476), .Y(N281) );
  AOI211X1TF U716 ( .A0(Y_IN[3]), .A1(N454), .B0(N279), .C0(N278), .Y(N282) );
  AOI211X1TF U717 ( .A0(X_IN[4]), .A1(N746), .B0(N114), .C0(N754), .Y(N278) );
  OAI32X1TF U718 ( .A0(N277), .A1(X_IN[2]), .A2(N324), .B0(X_IN[1]), .B1(N277), 
        .Y(N279) );
  OAI211X1TF U719 ( .A0(Y_IN[3]), .A1(N454), .B0(N276), .C0(N326), .Y(N277) );
  AOI22X1TF U720 ( .A0(N114), .A1(N754), .B0(X_IN[2]), .B1(N325), .Y(N276) );
  INVX2TF U721 ( .A(X_IN[4]), .Y(N454) );
  INVX2TF U722 ( .A(X_IN[6]), .Y(N476) );
  INVX2TF U723 ( .A(X_IN[8]), .Y(N502) );
  NOR2X1TF U724 ( .A(Y_IN[9]), .B(N515), .Y(N289) );
  INVX2TF U725 ( .A(X_IN[10]), .Y(N515) );
  NOR2X1TF U726 ( .A(Y_IN[11]), .B(N315), .Y(N295) );
  INVX2TF U727 ( .A(X_IN[12]), .Y(N315) );
  INVX2TF U728 ( .A(N349), .Y(N396) );
  OAI211X1TF U729 ( .A0(N873), .A1(N872), .B0(N871), .C0(N870), .Y(N678) );
  AOI32X1TF U730 ( .A0(N954), .A1(OPER_B[4]), .A2(N869), .B0(N901), .B1(
        OPER_B[4]), .Y(N870) );
  AOI211X1TF U731 ( .A0(N875), .A1(OPER_B[5]), .B0(N868), .C0(N867), .Y(N871)
         );
  OAI31X1TF U732 ( .A0(N951), .A1(OPER_A[4]), .A2(N866), .B0(N217), .Y(N867)
         );
  AOI21X1TF U733 ( .A0(N138), .A1(C152_DATA4_4), .B0(N219), .Y(N217) );
  NOR3X1TF U734 ( .A(OPER_B[4]), .B(N869), .C(N141), .Y(N868) );
  AOI21X1TF U735 ( .A0(N948), .A1(N866), .B0(N865), .Y(N872) );
  INVX2TF U736 ( .A(N949), .Y(N865) );
  AOI211X1TF U737 ( .A0(N139), .A1(C152_DATA4_5), .B0(N877), .C0(N223), .Y(
        N224) );
  OAI31X1TF U738 ( .A0(OPER_B[5]), .A1(N876), .A2(N141), .B0(N922), .Y(N877)
         );
  OAI211X1TF U739 ( .A0(SIGN_Y), .A1(N982), .B0(N233), .C0(N989), .Y(N922) );
  AOI22X1TF U740 ( .A0(N875), .A1(OPER_B[6]), .B0(N874), .B1(N879), .Y(N884)
         );
  NOR2X1TF U741 ( .A(N951), .B(OPER_A[5]), .Y(N874) );
  INVX2TF U742 ( .A(N911), .Y(N875) );
  AOI22X1TF U743 ( .A0(OPER_B[5]), .A1(N881), .B0(OPER_A[5]), .B1(N880), .Y(
        N883) );
  OAI21X1TF U744 ( .A0(N951), .A1(N879), .B0(N949), .Y(N880) );
  OAI21X1TF U745 ( .A0(N141), .A1(N878), .B0(N952), .Y(N881) );
  OAI211X1TF U746 ( .A0(N911), .A1(N185), .B0(N910), .C0(N909), .Y(N675) );
  AOI211X1TF U747 ( .A0(OPER_A[7]), .A1(N907), .B0(N906), .C0(N905), .Y(N910)
         );
  INVX2TF U748 ( .A(N220), .Y(N905) );
  AOI211X1TF U749 ( .A0(N138), .A1(C152_DATA4_7), .B0(N219), .C0(N218), .Y(
        N220) );
  NOR3X1TF U750 ( .A(N140), .B(OPER_B[7]), .C(N904), .Y(N218) );
  OR2X2TF U751 ( .A(N947), .B(N903), .Y(N219) );
  NOR2X1TF U752 ( .A(N984), .B(N847), .Y(N887) );
  INVX2TF U753 ( .A(N902), .Y(N906) );
  AOI32X1TF U754 ( .A0(OPER_B[7]), .A1(N954), .A2(N904), .B0(N901), .B1(
        OPER_B[7]), .Y(N902) );
  INVX2TF U755 ( .A(N952), .Y(N901) );
  OAI21X1TF U756 ( .A0(N951), .A1(N908), .B0(N949), .Y(N907) );
  NOR3X1TF U757 ( .A(N130), .B(N192), .C(N982), .Y(N981) );
  OAI22X1TF U758 ( .A0(N152), .A1(N214), .B0(N143), .B1(OFFSET[2]), .Y(C2_Z_4)
         );
  INVX2TF U759 ( .A(Y_IN[4]), .Y(N214) );
  OAI22X1TF U760 ( .A0(N152), .A1(N213), .B0(N143), .B1(OFFSET[3]), .Y(C2_Z_5)
         );
  OAI22X1TF U761 ( .A0(N152), .A1(N212), .B0(N143), .B1(OFFSET[4]), .Y(C2_Z_6)
         );
  OAI22X1TF U762 ( .A0(N151), .A1(N207), .B0(N143), .B1(OFFSET[5]), .Y(C2_Z_7)
         );
  OAI22X1TF U763 ( .A0(N152), .A1(N778), .B0(N143), .B1(OFFSET[6]), .Y(C2_Z_8)
         );
  OAI22X1TF U764 ( .A0(N151), .A1(N800), .B0(N143), .B1(OFFSET[7]), .Y(C2_Z_9)
         );
  OAI22X1TF U765 ( .A0(N152), .A1(N563), .B0(N143), .B1(OFFSET[8]), .Y(C2_Z_10) );
  OAI22X1TF U766 ( .A0(N152), .A1(N821), .B0(N143), .B1(OFFSET[9]), .Y(C2_Z_11) );
  INVX2TF U767 ( .A(Y_IN[11]), .Y(N821) );
  NOR2X1TF U768 ( .A(OPER_B[9]), .B(N925), .Y(N940) );
  NOR2X1TF U769 ( .A(N886), .B(OPER_B[6]), .Y(N904) );
  INVX2TF U770 ( .A(N890), .Y(N886) );
  NOR2X1TF U771 ( .A(OPER_B[5]), .B(N878), .Y(N890) );
  NOR2X1TF U772 ( .A(OPER_B[3]), .B(N858), .Y(N869) );
  AOI211X1TF U773 ( .A0(N131), .A1(N982), .B0(SIGN_Y), .C0(N927), .Y(N947) );
  NOR2X1TF U774 ( .A(OPER_A[9]), .B(N926), .Y(N934) );
  NOR2X1TF U775 ( .A(OPER_A[7]), .B(N908), .Y(N915) );
  NOR2X1TF U776 ( .A(OPER_A[5]), .B(N879), .Y(N893) );
  NOR2X1TF U777 ( .A(OPER_A[3]), .B(N857), .Y(N866) );
  OAI21X1TF U778 ( .A0(N536), .A1(N137), .B0(N260), .Y(OPER_A[4]) );
  OAI21X1TF U779 ( .A0(N455), .A1(N137), .B0(N261), .Y(OPER_A[5]) );
  OAI21X1TF U780 ( .A0(N541), .A1(N137), .B0(N262), .Y(OPER_A[6]) );
  OAI21X1TF U781 ( .A0(N477), .A1(N137), .B0(N263), .Y(OPER_A[7]) );
  OAI21X1TF U782 ( .A0(N175), .A1(N137), .B0(N264), .Y(OPER_A[8]) );
  OAI21X1TF U783 ( .A0(N137), .A1(N544), .B0(N265), .Y(OPER_A[9]) );
  OAI21X1TF U784 ( .A0(N137), .A1(N176), .B0(N266), .Y(OPER_A[10]) );
  OAI21X1TF U785 ( .A0(N137), .A1(N169), .B0(N267), .Y(OPER_A[11]) );
  OAI211X1TF U786 ( .A0(N191), .A1(N955), .B0(N864), .C0(N863), .Y(N679) );
  AOI211X1TF U787 ( .A0(OPER_A[3]), .A1(N862), .B0(N861), .C0(N860), .Y(N863)
         );
  OAI31X1TF U788 ( .A0(N951), .A1(OPER_A[3]), .A2(N859), .B0(N216), .Y(N860)
         );
  AOI21X1TF U789 ( .A0(C152_DATA4_3), .A1(N138), .B0(N923), .Y(N216) );
  OAI21X1TF U790 ( .A0(N152), .A1(N324), .B0(N142), .Y(C2_Z_1) );
  OAI22X1TF U791 ( .A0(N152), .A1(N746), .B0(N142), .B1(OFFSET[1]), .Y(C2_Z_3)
         );
  INVX2TF U792 ( .A(Y_IN[3]), .Y(N746) );
  OAI32X1TF U793 ( .A0(N197), .A1(N140), .A2(N858), .B0(N952), .B1(N197), .Y(
        N861) );
  INVX2TF U794 ( .A(N885), .Y(N938) );
  AOI32X1TF U795 ( .A0(N621), .A1(N357), .A2(N840), .B0(N963), .B1(N356), .Y(
        N885) );
  INVX2TF U796 ( .A(N957), .Y(N963) );
  OAI21X1TF U797 ( .A0(N951), .A1(N857), .B0(N949), .Y(N862) );
  INVX2TF U798 ( .A(N848), .Y(N929) );
  AOI21X1TF U799 ( .A0(N580), .A1(N356), .B0(N579), .Y(N848) );
  INVX2TF U800 ( .A(N859), .Y(N857) );
  NOR3X1TF U801 ( .A(OPER_A[2]), .B(OPER_A[1]), .C(OPER_A[0]), .Y(N859) );
  OAI21X1TF U802 ( .A0(N167), .A1(N136), .B0(N258), .Y(OPER_A[2]) );
  INVX2TF U803 ( .A(N948), .Y(N951) );
  NOR2X2TF U804 ( .A(N941), .B(N933), .Y(N948) );
  INVX2TF U805 ( .A(N921), .Y(N941) );
  OAI21X1TF U806 ( .A0(N168), .A1(N136), .B0(N259), .Y(OPER_A[3]) );
  AOI31X1TF U807 ( .A0(N954), .A1(N197), .A2(N858), .B0(N899), .Y(N864) );
  OAI21X1TF U808 ( .A0(N992), .A1(N927), .B0(N854), .Y(N899) );
  INVX2TF U809 ( .A(N927), .Y(N233) );
  INVX2TF U810 ( .A(N355), .Y(N976) );
  INVX2TF U811 ( .A(N581), .Y(N966) );
  NOR2X1TF U812 ( .A(OPER_B[1]), .B(OPER_B[0]), .Y(N850) );
  AOI22X1TF U813 ( .A0(N130), .A1(DIVISION_HEAD[3]), .B0(XTEMP[12]), .B1(N131), 
        .Y(N356) );
  INVX2TF U814 ( .A(N621), .Y(N839) );
  NOR2X2TF U815 ( .A(N619), .B(N647), .Y(N840) );
  AOI221X1TF U816 ( .A0(N128), .A1(N183), .B0(N195), .B1(N91), .C0(N835), .Y(
        N836) );
  AOI22X1TF U817 ( .A0(\INDEX[2] ), .A1(N90), .B0(N124), .B1(\RSHT_BITS[3] ), 
        .Y(N834) );
  AOI32X1TF U818 ( .A0(N957), .A1(N970), .A2(N380), .B0(N972), .B1(N970), .Y(
        N353) );
  OR2X2TF U819 ( .A(N647), .B(N177), .Y(N380) );
  INVX2TF U820 ( .A(N619), .Y(N728) );
  OAI21X1TF U821 ( .A0(N355), .A1(N956), .B0(N351), .Y(N623) );
  OAI21X1TF U822 ( .A0(N586), .A1(N580), .B0(N352), .Y(N351) );
  NOR2X2TF U823 ( .A(\RSHT_BITS[3] ), .B(N607), .Y(N621) );
  NOR3X1TF U824 ( .A(N121), .B(N122), .C(N971), .Y(N838) );
  NOR2X1TF U825 ( .A(SIGN_Y), .B(N61), .Y(N924) );
  INVX2TF U826 ( .A(N322), .Y(N643) );
  OAI22X1TF U827 ( .A0(Y_IN[12]), .A1(N175), .B0(N347), .B1(N346), .Y(N348) );
  OAI31X1TF U828 ( .A0(N345), .A1(DIVISION_HEAD[10]), .A2(N563), .B0(N344), 
        .Y(N346) );
  AOI22X1TF U829 ( .A0(Y_IN[11]), .A1(N477), .B0(N343), .B1(N342), .Y(N344) );
  OAI22X1TF U830 ( .A0(DIVISION_HEAD[8]), .A1(N778), .B0(DIVISION_HEAD[9]), 
        .B1(N800), .Y(N342) );
  INVX2TF U831 ( .A(N341), .Y(N343) );
  NOR2X1TF U832 ( .A(Y_IN[11]), .B(N477), .Y(N345) );
  AOI211X1TF U833 ( .A0(DIVISION_HEAD[8]), .A1(N778), .B0(N340), .C0(N341), 
        .Y(N347) );
  OAI21X1TF U834 ( .A0(Y_IN[11]), .A1(N477), .B0(N339), .Y(N341) );
  INVX2TF U835 ( .A(Y_IN[9]), .Y(N800) );
  INVX2TF U836 ( .A(Y_IN[10]), .Y(N563) );
  AOI21X1TF U837 ( .A0(N113), .A1(N168), .B0(N338), .Y(N340) );
  AOI211X1TF U838 ( .A0(N337), .A1(DIVISION_HEAD[6]), .B0(N336), .C0(N335), 
        .Y(N338) );
  NOR2X1TF U839 ( .A(N113), .B(N168), .Y(N336) );
  AOI211X1TF U840 ( .A0(N333), .A1(DIVISION_HEAD[4]), .B0(N332), .C0(N331), 
        .Y(N334) );
  NOR2X1TF U841 ( .A(Y_IN[5]), .B(N527), .Y(N332) );
  AOI21X1TF U842 ( .A0(Y_IN[3]), .A1(N734), .B0(N330), .Y(N333) );
  OAI32X1TF U843 ( .A0(N329), .A1(DIVISION_HEAD[2]), .A2(N754), .B0(N328), 
        .B1(N329), .Y(N330) );
  OAI211X1TF U844 ( .A0(Y_IN[2]), .A1(N829), .B0(N327), .C0(N326), .Y(N328) );
  INVX2TF U845 ( .A(Y_IN[0]), .Y(N742) );
  INVX2TF U846 ( .A(Y_IN[1]), .Y(N324) );
  INVX2TF U847 ( .A(Y_IN[2]), .Y(N754) );
  INVX2TF U848 ( .A(Y_IN[8]), .Y(N778) );
  INVX2TF U849 ( .A(Y_IN[12]), .Y(N564) );
  NOR2X1TF U850 ( .A(N254), .B(N368), .Y(FOUT[12]) );
  AND2X2TF U851 ( .A(ZTEMP[12]), .B(N159), .Y(POUT[12]) );
  OAI21X1TF U852 ( .A0(N167), .A1(N254), .B0(N239), .Y(FOUT[2]) );
  AOI21X1TF U853 ( .A0(N232), .A1(DIVISION_REMA[2]), .B0(N238), .Y(N239) );
  OAI22X1TF U854 ( .A0(N536), .A1(N110), .B0(N173), .B1(N107), .Y(N238) );
  AND2X2TF U855 ( .A(ZTEMP[2]), .B(N204), .Y(POUT[2]) );
  AND2X2TF U856 ( .A(ZTEMP[10]), .B(N159), .Y(POUT[10]) );
  OAI21X1TF U857 ( .A0(N168), .A1(N254), .B0(N241), .Y(FOUT[3]) );
  AOI21X1TF U858 ( .A0(N232), .A1(DIVISION_REMA[3]), .B0(N240), .Y(N241) );
  OAI22X1TF U859 ( .A0(N455), .A1(N109), .B0(N170), .B1(N107), .Y(N240) );
  AND2X2TF U860 ( .A(ZTEMP[3]), .B(N204), .Y(POUT[3]) );
  AND2X2TF U861 ( .A(ZTEMP[9]), .B(N159), .Y(POUT[9]) );
  NOR2X1TF U862 ( .A(N254), .B(N169), .Y(FOUT[11]) );
  AND2X2TF U863 ( .A(ZTEMP[11]), .B(N159), .Y(POUT[11]) );
  OAI21X1TF U864 ( .A0(N175), .A1(N254), .B0(N251), .Y(FOUT[8]) );
  AOI21X1TF U865 ( .A0(N232), .A1(DIVISION_REMA[8]), .B0(N250), .Y(N251) );
  OAI22X1TF U866 ( .A0(N165), .A1(N108), .B0(N176), .B1(N109), .Y(N250) );
  AND2X2TF U867 ( .A(ZTEMP[8]), .B(N159), .Y(POUT[8]) );
  OAI21X1TF U868 ( .A0(N527), .A1(N254), .B0(N237), .Y(FOUT[1]) );
  AOI21X1TF U869 ( .A0(N232), .A1(DIVISION_REMA[1]), .B0(N236), .Y(N237) );
  OAI22X1TF U870 ( .A0(N168), .A1(N109), .B0(N752), .B1(N107), .Y(N236) );
  AND2X2TF U871 ( .A(ZTEMP[1]), .B(N204), .Y(POUT[1]) );
  OAI21X1TF U872 ( .A0(N455), .A1(N254), .B0(N245), .Y(FOUT[5]) );
  AOI21X1TF U873 ( .A0(N232), .A1(DIVISION_REMA[5]), .B0(N244), .Y(N245) );
  OAI22X1TF U874 ( .A0(N477), .A1(N109), .B0(N171), .B1(N107), .Y(N244) );
  OAI21X1TF U875 ( .A0(N536), .A1(N157), .B0(N243), .Y(FOUT[4]) );
  AOI21X1TF U876 ( .A0(N232), .A1(DIVISION_REMA[4]), .B0(N242), .Y(N243) );
  OAI22X1TF U877 ( .A0(N541), .A1(N110), .B0(N174), .B1(N107), .Y(N242) );
  AND2X2TF U878 ( .A(ZTEMP[4]), .B(N204), .Y(POUT[4]) );
  OAI21X1TF U879 ( .A0(N477), .A1(N254), .B0(N249), .Y(FOUT[7]) );
  AOI21X1TF U880 ( .A0(N232), .A1(DIVISION_REMA[7]), .B0(N248), .Y(N249) );
  OAI22X1TF U881 ( .A0(N172), .A1(N108), .B0(N544), .B1(N109), .Y(N248) );
  AND2X2TF U882 ( .A(ZTEMP[7]), .B(N204), .Y(POUT[7]) );
  OAI21X1TF U883 ( .A0(N541), .A1(N157), .B0(N247), .Y(FOUT[6]) );
  AOI21X1TF U884 ( .A0(N232), .A1(DIVISION_REMA[6]), .B0(N246), .Y(N247) );
  OAI22X1TF U885 ( .A0(N175), .A1(N110), .B0(N164), .B1(N108), .Y(N246) );
  INVX2TF U886 ( .A(N272), .Y(N254) );
  NOR2X1TF U887 ( .A(N349), .B(N381), .Y(ALU_IS_DONE) );
  OAI211X1TF U888 ( .A0(N167), .A1(N110), .B0(N235), .C0(N234), .Y(FOUT[0]) );
  AND2X2TF U889 ( .A(ZTEMP[0]), .B(N159), .Y(POUT[0]) );
  AOI22X1TF U890 ( .A0(N149), .A1(\INTADD_0_SUM[5] ), .B0(N816), .B1(
        SUM_AB[10]), .Y(N461) );
  AOI21X1TF U891 ( .A0(N149), .A1(N486), .B0(N485), .Y(N487) );
  AOI22X1TF U892 ( .A0(N148), .A1(N479), .B0(SUM_AB[8]), .B1(N153), .Y(N481)
         );
  AOI31X1TF U893 ( .A0(X_IN[0]), .A1(N149), .A2(N179), .B0(N402), .Y(N403) );
  AOI22X1TF U894 ( .A0(N149), .A1(\INTADD_0_SUM[1] ), .B0(SUM_AB[2]), .B1(N154), .Y(N424) );
  AOI22X1TF U895 ( .A0(N149), .A1(\INTADD_0_SUM[3] ), .B0(SUM_AB[4]), .B1(N154), .Y(N443) );
  AOI22X1TF U896 ( .A0(N149), .A1(\INTADD_0_SUM[6] ), .B0(SUM_AB[7]), .B1(N154), .Y(N474) );
  AOI22X1TF U897 ( .A0(N149), .A1(\INTADD_0_SUM[0] ), .B0(SUM_AB[1]), .B1(N154), .Y(N414) );
  AOI22X1TF U898 ( .A0(N148), .A1(\INTADD_0_SUM[4] ), .B0(SUM_AB[5]), .B1(N153), .Y(N450) );
  AOI31X1TF U899 ( .A0(N148), .A1(N176), .A2(N508), .B0(N503), .Y(N504) );
  AOI22X1TF U900 ( .A0(N149), .A1(\INTADD_0_SUM[2] ), .B0(SUM_AB[3]), .B1(N154), .Y(N434) );
  AOI31X1TF U901 ( .A0(N149), .A1(N169), .A2(N523), .B0(N521), .Y(N525) );
  AOI21X1TF U902 ( .A0(N149), .A1(N367), .B0(N526), .Y(N369) );
  NAND3X1TF U903 ( .A(N922), .B(N227), .C(N226), .Y(N674) );
  NAND4BX1TF U904 ( .AN(N855), .B(N222), .C(N856), .D(N221), .Y(N680) );
  AOI2BB2X1TF U905 ( .B0(N139), .B1(C152_DATA4_2), .A0N(N181), .A1N(N946), .Y(
        N221) );
  OAI2BB1X1TF U906 ( .A0N(N139), .A1N(C152_DATA4_10), .B0(N228), .Y(N672) );
  NAND3X1TF U907 ( .A(N883), .B(N884), .C(N224), .Y(N677) );
  NAND2BX1TF U908 ( .AN(DP_OP_333_124_4748_N57), .B(N151), .Y(N215) );
  OAI2BB2XLTF U909 ( .B0(OFFSET[0]), .B1(N142), .A0N(Y_IN[2]), .A1N(N988), .Y(
        C2_Z_2) );
  INVX2TF U910 ( .A(N977), .Y(N984) );
  AOI2BB2X1TF U911 ( .B0(N232), .B1(DIVISION_REMA[0]), .A0N(N180), .A1N(N108), 
        .Y(N235) );
  OAI222X1TF U912 ( .A0(N110), .A1(N368), .B0(N108), .B1(N734), .C0(N254), 
        .C1(N176), .Y(FOUT[10]) );
  OAI222X1TF U913 ( .A0(N254), .A1(N544), .B0(N108), .B1(N829), .C0(N169), 
        .C1(N110), .Y(FOUT[9]) );
  NAND2X1TF U914 ( .A(N177), .B(N188), .Y(N381) );
  NAND3X1TF U915 ( .A(STEP[2]), .B(STEP[3]), .C(N728), .Y(N957) );
  NAND3X1TF U916 ( .A(N561), .B(N398), .C(N650), .Y(N733) );
  NOR4XLTF U917 ( .A(N779), .B(N633), .C(N818), .D(N733), .Y(N275) );
  AOI222XLTF U918 ( .A0(STEP[2]), .A1(N178), .B0(N121), .B1(N188), .C0(N166), 
        .C1(N122), .Y(N273) );
  NAND3X1TF U919 ( .A(N275), .B(N372), .C(N649), .Y(N635) );
  NAND2X1TF U920 ( .A(Y_IN[1]), .B(Y_IN[0]), .Y(N325) );
  AOI2BB1X1TF U921 ( .A0N(X_IN[5]), .A1N(N282), .B0(Y_IN[4]), .Y(N280) );
  AOI2BB1X1TF U922 ( .A0N(X_IN[7]), .A1N(N286), .B0(Y_IN[6]), .Y(N284) );
  NAND2X1TF U923 ( .A(MODE_TYPE[0]), .B(N323), .Y(N780) );
  AO22X1TF U924 ( .A0(X_IN[4]), .A1(N754), .B0(N114), .B1(N325), .Y(N297) );
  NAND2X1TF U925 ( .A(N127), .B(N746), .Y(N299) );
  AOI2BB1X1TF U926 ( .A0N(N303), .A1N(X_IN[6]), .B0(Y_IN[4]), .Y(N301) );
  AOI2BB1X1TF U927 ( .A0N(N307), .A1N(X_IN[8]), .B0(Y_IN[6]), .Y(N305) );
  NAND2X1TF U928 ( .A(N182), .B(N195), .Y(N632) );
  NAND2X1TF U929 ( .A(N850), .B(N181), .Y(N858) );
  NAND2X1TF U930 ( .A(N869), .B(N191), .Y(N878) );
  NOR2BX1TF U931 ( .AN(N904), .B(OPER_B[7]), .Y(N912) );
  NAND2X1TF U932 ( .A(N912), .B(N185), .Y(N925) );
  NAND2X1TF U933 ( .A(N940), .B(N186), .Y(N953) );
  NAND2X1TF U934 ( .A(N924), .B(N74), .Y(N975) );
  NAND2X1TF U935 ( .A(N581), .B(N975), .Y(N956) );
  NAND2X1TF U936 ( .A(N984), .B(N389), .Y(N589) );
  NAND3X1TF U937 ( .A(N92), .B(N91), .C(N90), .Y(N607) );
  NOR2BX1TF U938 ( .AN(N589), .B(N621), .Y(N586) );
  NAND2X1TF U939 ( .A(PRE_WORK), .B(N361), .Y(N970) );
  NAND2X1TF U940 ( .A(N621), .B(N840), .Y(N354) );
  NAND2X1TF U941 ( .A(N231), .B(N976), .Y(N374) );
  NAND3X1TF U942 ( .A(SIGN_Y), .B(N74), .C(N923), .Y(N841) );
  NAND2X1TF U943 ( .A(N873), .B(N866), .Y(N879) );
  NAND2X1TF U944 ( .A(N892), .B(N893), .Y(N908) );
  NAND2X1TF U945 ( .A(N914), .B(N915), .Y(N926) );
  NAND2X1TF U946 ( .A(N932), .B(N934), .Y(N950) );
  NAND3X1TF U947 ( .A(N621), .B(N618), .C(N187), .Y(N616) );
  NAND2X1TF U948 ( .A(N427), .B(N426), .Y(N435) );
  NAND2X1TF U949 ( .A(N445), .B(N444), .Y(N456) );
  NAND2X1TF U950 ( .A(N466), .B(N465), .Y(N475) );
  NAND2X1TF U951 ( .A(N513), .B(N512), .Y(N1031) );
  AOI222XLTF U952 ( .A0(XTEMP[11]), .A1(X_IN[11]), .B0(XTEMP[11]), .B1(N511), 
        .C0(X_IN[11]), .C1(N511), .Y(N362) );
  XOR2X1TF U953 ( .A(X_IN[12]), .B(N362), .Y(N367) );
  NAND3X1TF U954 ( .A(N582), .B(POST_WORK), .C(N618), .Y(N384) );
  NAND3BX1TF U955 ( .AN(N374), .B(N966), .C(N984), .Y(N614) );
  NAND3X1TF U956 ( .A(N625), .B(N375), .C(N614), .Y(N960) );
  NAND2X1TF U957 ( .A(N145), .B(N406), .Y(N393) );
  NAND3X1TF U958 ( .A(N396), .B(N122), .C(DP_OP_333_124_4748_N57), .Y(N654) );
  NOR2BX1TF U959 ( .AN(N650), .B(N961), .Y(N558) );
  NAND3X1TF U960 ( .A(N558), .B(N388), .C(N387), .Y(N392) );
  NAND4X1TF U961 ( .A(N439), .B(N438), .C(N437), .D(N436), .Y(N440) );
  NAND4X1TF U962 ( .A(N450), .B(N449), .C(N448), .D(N447), .Y(N451) );
  NAND4X1TF U963 ( .A(N461), .B(N460), .C(N459), .D(N458), .Y(N462) );
  OAI2BB1X1TF U964 ( .A0N(DIVISION_HEAD[10]), .A1N(N485), .B0(N464), .Y(N713)
         );
  AOI2BB2X1TF U965 ( .B0(X_IN[9]), .B1(N492), .A0N(N492), .A1N(X_IN[9]), .Y(
        N497) );
  NAND3X1TF U966 ( .A(N148), .B(N544), .C(N497), .Y(N493) );
  AOI2BB1X1TF U967 ( .A0N(N522), .A1N(N497), .B0(N526), .Y(N498) );
  AOI2BB2X1TF U968 ( .B0(N501), .B1(N515), .A0N(N515), .A1N(N501), .Y(N508) );
  AOI2BB1X1TF U969 ( .A0N(N522), .A1N(N508), .B0(N526), .Y(N509) );
  AOI2BB2X1TF U970 ( .B0(N105), .B1(N511), .A0N(N511), .A1N(N105), .Y(N523) );
  OAI2BB2XLTF U971 ( .B0(N515), .B1(N624), .A0N(XTEMP[12]), .A1N(N115), .Y(
        N516) );
  AOI2BB1X1TF U972 ( .A0N(N522), .A1N(N523), .B0(N526), .Y(N524) );
  AOI2BB1X1TF U973 ( .A0N(DIVISION_REMA[2]), .A1N(N531), .B0(DIVISION_HEAD[6]), 
        .Y(N529) );
  OA21XLTF U974 ( .A0(N536), .A1(DIVISION_REMA[4]), .B0(N533), .Y(N535) );
  OA21XLTF U975 ( .A0(N541), .A1(DIVISION_REMA[6]), .B0(N538), .Y(N540) );
  OA21XLTF U976 ( .A0(XTEMP[12]), .A1(N551), .B0(N734), .Y(N550) );
  NAND4X1TF U977 ( .A(N561), .B(N560), .C(N654), .D(N559), .Y(N572) );
  NAND3X1TF U978 ( .A(N567), .B(N566), .C(N565), .Y(N568) );
  NAND3X1TF U979 ( .A(N773), .B(N575), .C(N574), .Y(N576) );
  NAND3X1TF U980 ( .A(N582), .B(N618), .C(N839), .Y(N588) );
  NAND4X1TF U981 ( .A(N584), .B(N583), .C(N655), .D(N588), .Y(N585) );
  NAND2X1TF U982 ( .A(N194), .B(N183), .Y(N606) );
  NOR4XLTF U983 ( .A(\RSHT_BITS[3] ), .B(N90), .C(N630), .D(N606), .Y(N587) );
  NAND2X1TF U984 ( .A(N595), .B(N605), .Y(N602) );
  NAND2X1TF U985 ( .A(N92), .B(N91), .Y(N604) );
  AOI2BB2X1TF U986 ( .B0(N612), .B1(N183), .A0N(N606), .A1N(N608), .Y(N600) );
  NAND4X1TF U987 ( .A(N120), .B(N650), .C(N649), .D(N648), .Y(N651) );
  NAND4X1TF U988 ( .A(N656), .B(N655), .C(N654), .D(N729), .Y(N697) );
  NAND3X1TF U989 ( .A(N773), .B(N738), .C(N737), .Y(N739) );
  AO22X1TF U990 ( .A0(DIVISION_REMA[4]), .A1(N751), .B0(N206), .B1(N807), .Y(
        N760) );
  AOI2BB1X1TF U991 ( .A0N(X_IN[1]), .A1N(N781), .B0(N780), .Y(N784) );
  NAND4X1TF U992 ( .A(N811), .B(N810), .C(N809), .D(N808), .Y(N812) );
  OAI221XLTF U993 ( .A0(\INDEX[2] ), .A1(N90), .B0(N124), .B1(\RSHT_BITS[3] ), 
        .C0(N834), .Y(N835) );
  OAI221XLTF U994 ( .A0(N129), .A1(N194), .B0(N182), .B1(N92), .C0(N836), .Y(
        N847) );
  NAND2X1TF U995 ( .A(N921), .B(N887), .Y(N882) );
  NAND2BX1TF U996 ( .AN(N837), .B(N882), .Y(N903) );
  NAND2X1TF U997 ( .A(N846), .B(N984), .Y(N888) );
  NAND3X1TF U998 ( .A(SIGN_Y), .B(N74), .C(N233), .Y(N854) );
  OAI2BB1X1TF U999 ( .A0N(N977), .A1N(N847), .B0(N846), .Y(N937) );
  NAND3X1TF U1000 ( .A(N74), .B(N192), .C(N131), .Y(N992) );
  NAND4X1TF U1001 ( .A(N233), .B(N192), .C(N131), .D(N982), .Y(N856) );
  NAND2X1TF U1002 ( .A(N921), .B(N937), .Y(N955) );
  NAND3BX1TF U1003 ( .AN(OPER_A[7]), .B(N948), .C(N908), .Y(N909) );
  NAND2X1TF U1004 ( .A(N103), .B(N963), .Y(N964) );
  NAND2X1TF U1005 ( .A(N996), .B(N995), .Y(N668) );
  NAND2X1TF U1006 ( .A(N999), .B(N998), .Y(N667) );
  NAND2X1TF U1007 ( .A(SUM_AB[3]), .B(N112), .Y(N1000) );
  NAND2X1TF U1008 ( .A(N1005), .B(N1004), .Y(N665) );
  NAND2X1TF U1009 ( .A(SUM_AB[5]), .B(N112), .Y(N1006) );
  NAND2X1TF U1010 ( .A(N1011), .B(N1010), .Y(N663) );
  NAND2X1TF U1011 ( .A(SUM_AB[7]), .B(N112), .Y(N1012) );
  NAND2X1TF U1012 ( .A(N1017), .B(N1016), .Y(N661) );
  NAND2X1TF U1013 ( .A(SUM_AB[9]), .B(N112), .Y(N1018) );
  NAND2X1TF U1014 ( .A(N1023), .B(N1022), .Y(N659) );
  NAND2X1TF U1015 ( .A(SUM_AB[11]), .B(N112), .Y(N1024) );
endmodule


module SERIAL_CPU_8BIT_VG ( CLK, ENABLE, RST_N, START, I_DATAIN, D_DATAIN, 
        IS_I_ADDR, NXT, I_ADDR, D_ADDR, D_WE, D_DATAOUT, IO_STATUS, IO_CONTROL, 
        IO_DATAINA, IO_DATAINB, IO_DATAOUTA, IO_DATAOUTB, IO_OFFSET );
  input [7:0] I_DATAIN;
  input [7:0] D_DATAIN;
  output [1:0] NXT;
  output [8:0] I_ADDR;
  output [8:0] D_ADDR;
  output [7:0] D_DATAOUT;
  input [15:0] IO_STATUS;
  output [15:0] IO_CONTROL;
  input [15:0] IO_DATAINA;
  input [15:0] IO_DATAINB;
  output [15:0] IO_DATAOUTA;
  output [15:0] IO_DATAOUTB;
  output [15:0] IO_OFFSET;
  input CLK, ENABLE, RST_N, START;
  output IS_I_ADDR, D_WE;
  wire   \OPER1_R1[2] , N114, N162, N163, N164, CF_BUF, N466, N467, N468, N469,
         N470, N471, N472, N473, N474, N475, N476, N477, N478, N479, N480,
         N481, N482, N500, N501, N502, N503, N504, N505, N506, N507, N508,
         N509, N510, N511, N512, N513, N514, N515, N516, N584, N585, ZF, NF,
         CF, N612, N412, N414, N415, N416, N417, N418, N420, N421, N423, N424,
         N429, N431, N432, N442, N443, N444, N445, N446, N447, N448, N449,
         N450, N451, N452, N453, N454, N455, N456, N457, N458, N460, N461,
         N462, N463, N464, N465, N4660, N4670, N4680, N4690, N4700, N4710,
         N4720, N4730, N4740, N4750, N4760, N4770, N4780, N4790, N4800, N4810,
         N4820, N483, N484, N485, N486, N487, N488, N492, N493, N494, N495,
         N496, N497, N498, N499, N5030, N5040, N5060, N5070, N5090, N5100,
         N5120, N5130, N5150, N5160, N518, N519, N521, N522, N524, N525, N527,
         N528, N530, N531, N533, N534, N536, N537, N539, N540, N542, N543,
         N545, N558, N562, N564, N579, N582, N605, N606, N607, N608, N609,
         N610, N611, N6120, N613, N614, N615, N616, N617, N618, N619, N620,
         N623, N624, N625, N626, N627, N628, N629, N630, N631, N632, N633,
         N634, N635, N636, N637, N638, N639, N640, N641, N642, N643, N644,
         N645, N646, N647, N648, N649, N650, N651, N652, N653, N654, N655,
         N656, N657, N658, N659, N660, N661, N662, N663, N664, N665, N666,
         N667, N668, N669, N670, N671, N672, N673, N674, N675, N676, N677,
         N678, N679, N680, N681, N682, N683, N684, N685, N686, N687, N688,
         N689, N690, N691, N692, N693, N694, N695, N696, N697, N698, N699,
         N700, N701, N702, N817, N821, N822, N823, N824, N825, N873, N874,
         N936, N937, N938, N939, N940, N941, N942, N943, N944, N945, N946,
         N947, N948, N949, N950, N951, N952, N953, N954, N955, N956, N957,
         N958, N959, N960, N961, N962, N963, N964, N965, N966, N967, N968,
         N969, N970, N971, N972, N973, N974, N975, N976, N977, N978, N979,
         N980, N981, N982, N983, N984, N985, N986, N987, N988, N989, N990,
         N991, N992, N993, N994, N995, N996, N997, N998, N999, N1000, N1001,
         N1002, N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011,
         N1012, N1013, N1014, N1015, N1016, SUB_X_283_4_N16, SUB_X_283_4_N15,
         SUB_X_283_4_N14, SUB_X_283_4_N13, SUB_X_283_4_N12, SUB_X_283_4_N11,
         SUB_X_283_4_N10, SUB_X_283_4_N9, SUB_X_283_4_N8, SUB_X_283_4_N7,
         SUB_X_283_4_N6, SUB_X_283_4_N5, SUB_X_283_4_N4, SUB_X_283_4_N3,
         SUB_X_283_4_N2, SUB_X_283_4_N1, ADD_X_283_3_N16, ADD_X_283_3_N15,
         ADD_X_283_3_N14, ADD_X_283_3_N13, ADD_X_283_3_N12, ADD_X_283_3_N11,
         ADD_X_283_3_N10, ADD_X_283_3_N9, ADD_X_283_3_N8, ADD_X_283_3_N7,
         ADD_X_283_3_N6, ADD_X_283_3_N5, ADD_X_283_3_N4, ADD_X_283_3_N3,
         ADD_X_283_3_N2, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12,
         N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N158,
         N159, N160, N1620, N1630, N1640, N165, N166, N167, N168, N169, N170,
         N171, N172, N173, N174, N175, N176, N177, N178, N179, N180, N181,
         N182, N183, N184, N185, N186, N187, N188, N189, N190, N191, N192,
         N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204,
         N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215,
         N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226,
         N227, N228, N229, N230, N231, N239, N240, N241, N242, N243, N244,
         N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255,
         N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266,
         N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277,
         N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288,
         N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299,
         N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, N310,
         N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, N321,
         N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332,
         N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343,
         N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, N354,
         N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365,
         N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376,
         N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387,
         N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398,
         N399, N400, N401, N402, N403, N404, N405, N406, N407, N408, N409,
         N410, N411, N413, N419, N422, N425, N426, N427, N428, N430, N433,
         N434, N435, N436, N437, N438, N439, N440, N441, N459, N489, N490,
         N491, N5000, N5010, N5020, N5050, N5080, N5110, N5140, N517, N520,
         N523, N526, N529, N532, N535, N538, N541, N544, N546, N547, N548,
         N549, N550, N551, N552, N553, N554, N555, N556, N557, N559, N560,
         N561, N563, N565, N566, N567, N568, N569, N570, N571, N572, N573,
         N574, N575, N576, N577, N578, N580, N581, N583, N5840, N5850, N586,
         N587, N588, N589, N590, N591, N592, N593, N594, N595, N596, N597,
         N598, N599, N600, N601, N602, N603, N604, N621, N622, N703, N704,
         N705, N706, N707, N708, N709, N710, N711, N712, N713, N714, N715,
         N716, N717, N718, N719, N720, N721, N722, N723, N724, N725, N726,
         N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737,
         N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748,
         N749, N750, N751, N752, N753, N754, N755, N756, N757, N758, N759,
         N760, N761, N762, N763, N764, N765, N766, N767, N768, N769, N770,
         N771, N772, N773, N774, N775, N776, N777, N778, N779, N780, N781,
         N782, N783, N784, N785, N786, N787, N788, N789, N790, N791, N792,
         N793, N794, N795, N796, N797, N798, N799, N800, N801, N802, N803,
         N804, N805, N806, N807, N808, N809, N810, N811, N812, N813, N814,
         N815, N816, N818, N819, N820, N826, N827, N828, N829, N830, N831,
         N832, N833, N834, N835, N836, N837, N838, N839, N840, N841, N842,
         N843, N844, N845, N846, N847, N848, N849, N850, N851, N852, N853,
         N854, N855, N856, N857, N858, N859, N860, N861, N862, N863, N864,
         N865, N866, N867, N868, N869, N870, N871, N872, N875, N876, N877,
         N878, N879, N880, N881, N882, N883, N884, N885, N886, N887, N888,
         N889, N890, N891, N892, N893, N894, N895, N896, N897, N898, N899,
         N900, N901, N902, N903, N904, N905, N906, N907, N908, N909, N910,
         N911, N912, N913, N914, N915, N916, N917, N918, N919, N920, N921,
         N922, N923, N924, N925, N926, N927, N928, N929, N930, N931, N932,
         N933, N934, N935, N1017, N1018, N1019, N1020, N1021, N1022, N1023,
         N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1031, N1032, N1033,
         N1034, N1035, N1036, N1037, N1038, N1039, N1040, N1041, N1042, N1043,
         N1044, N1045, N1046, N1047, N1048, N1049, N1050, N1051, N1052, N1053,
         N1054, N1055, N1056, N1057, N1058, N1059, N1060, N1061, N1062, N1063,
         N1064, N1065, N1066, N1067, N1068, N1069, N1070, N1071, N1072, N1073,
         N1074, N1075, N1076, N1077, N1078, N1079, N1080, N1081, N1082, N1083,
         N1084, N1085, N1086, N1087, N1088, N1089, N1090, N1091, N1092, N1093,
         N1094, N1095, N1096, N1097, N1098, N1099, N1100, N1101, N1102, N1103,
         N1104, N1105, N1106, N1107, N1108, N1109, N1110, N1111, N1112, N1113,
         N1114, N1115, N1116, N1117, N1118, N1119, N1120, N1121, N1122, N1123,
         N1124, N1125, N1126, N1127, N1128, N1129, N1130, N1131, N1132, N1133,
         N1134, N1135, N1136, N1137, N1138, N1139, N1140, N1141, N1142, N1143,
         N1144, N1145, N1146, N1147, N1148, N1149, N1150, N1151, N1152, N1153,
         N1154, N1155, N1156, N1157, N1158, N1159, N1160, N1161, N1162, N1163,
         N1164, N1165, N1166, N1167, N1168, N1169, N1170, N1171, N1172, N1173,
         N1174, N1175, N1176, N1177, N1178, N1179, N1180, N1181, N1182, N1183,
         N1184, N1185, N1186, N1187, N1188, N1189, N1190, N1191, N1192, N1193,
         N1194, N1195, N1196, N1197, N1198, N1199, N1200, N1201, N1202, N1203,
         N1204, N1205, N1206, N1207, N1208, N1209, N1210, N1211, N1212, N1213,
         N1214, N1215, N1216;
  wire   [4:2] CODE_TYPE;
  wire   [2:0] OPER3_R3;
  wire   [1:0] STATE;
  wire   [2:0] NEXT_STATE;
  wire   [15:0] REG_A;
  wire   [15:0] REG_B;

  DFFRX4TF \reg_B_reg[0]  ( .D(N543), .CK(CLK), .RN(RST_N), .Q(REG_B[0]), .QN(
        N20) );
  DFFRX2TF \gr_reg[3][12]  ( .D(N946), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTB[12]), .QN(N642) );
  DFFSX2TF \pc_reg[2]  ( .D(N824), .CK(CLK), .SN(RST_N), .Q(N280), .QN(
        I_ADDR[3]) );
  DFFRX2TF \gr_reg[4][7]  ( .D(N975), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[7]), 
        .QN(N631) );
  DFFRX2TF \gr_reg[4][3]  ( .D(N979), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[3]), 
        .QN(N635) );
  DFFRX2TF \gr_reg[4][5]  ( .D(N977), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[5]), 
        .QN(N633) );
  DFFRX2TF \gr_reg[4][6]  ( .D(N976), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[6]), 
        .QN(N632) );
  DFFRX2TF \gr_reg[4][4]  ( .D(N978), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[4]), 
        .QN(N634) );
  DFFRX2TF \gr_reg[3][7]  ( .D(N983), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[7]), 
        .QN(N647) );
  DFFRX2TF \gr_reg[1][3]  ( .D(N1003), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[3]), 
        .QN(N683) );
  DFFRX2TF \gr_reg[3][4]  ( .D(N986), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[4]), 
        .QN(N650) );
  DFFRX2TF \gr_reg[3][15]  ( .D(N943), .CK(CLK), .RN(RST_N), .Q(N279), .QN(
        N639) );
  DFFRX2TF \gr_reg[3][14]  ( .D(N944), .CK(CLK), .RN(RST_N), .Q(N278), .QN(
        N640) );
  DFFRX2TF \gr_reg[3][11]  ( .D(N947), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTB[11]), .QN(N643) );
  DFFRX2TF \gr_reg[3][13]  ( .D(N945), .CK(CLK), .RN(RST_N), .Q(N277), .QN(
        N641) );
  DFFRX2TF \gr_reg[3][10]  ( .D(N948), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTB[10]), .QN(N644) );
  DFFRX2TF \gr_reg[3][9]  ( .D(N949), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[9]), 
        .QN(N645) );
  DFFRX2TF \gr_reg[3][6]  ( .D(N984), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[6]), 
        .QN(N648) );
  DFFRX2TF \gr_reg[3][8]  ( .D(N950), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[8]), 
        .QN(N646) );
  DFFRX2TF \gr_reg[3][0]  ( .D(N990), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[0]), 
        .QN(N654) );
  DFFRX2TF \gr_reg[3][1]  ( .D(N989), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[1]), 
        .QN(N653) );
  DFFRX2TF \gr_reg[3][2]  ( .D(N988), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[2]), 
        .QN(N652) );
  DFFSX2TF \pc_reg[7]  ( .D(N873), .CK(CLK), .SN(RST_N), .Q(N270), .QN(
        I_ADDR[8]) );
  DFFSX2TF \pc_reg[5]  ( .D(N821), .CK(CLK), .SN(RST_N), .Q(N269), .QN(
        I_ADDR[6]) );
  DFFSX2TF \pc_reg[3]  ( .D(N823), .CK(CLK), .SN(RST_N), .Q(N268), .QN(
        I_ADDR[4]) );
  DFFRX2TF \gr_reg[3][5]  ( .D(N985), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[5]), 
        .QN(N649) );
  DFFSX2TF \state_reg[3]  ( .D(N558), .CK(CLK), .SN(RST_N), .Q(N562), .QN(N263) );
  DFFRX2TF \id_ir_reg[1]  ( .D(N4720), .CK(CLK), .RN(RST_N), .Q(OPER3_R3[1]), 
        .QN(N260) );
  DFFRX2TF \id_ir_reg[15]  ( .D(N492), .CK(CLK), .RN(RST_N), .Q(CODE_TYPE[4]), 
        .QN(N242) );
  DFFRX2TF \id_ir_reg[11]  ( .D(N496), .CK(CLK), .RN(RST_N), .Q(N240), .QN(
        N579) );
  TLATXLTF cf_buf_reg ( .G(N584), .D(N585), .Q(CF_BUF) );
  TLATXLTF \nxt_reg[0]  ( .G(N162), .D(N163), .Q(NXT[0]) );
  TLATXLTF \nxt_reg[1]  ( .G(N162), .D(N164), .Q(NXT[1]) );
  DFFRX2TF \gr_reg[4][9]  ( .D(N941), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[9]), 
        .QN(N629) );
  DFFRX2TF \gr_reg[4][8]  ( .D(N942), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[8]), 
        .QN(N630) );
  DFFRX2TF \gr_reg[4][1]  ( .D(N981), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[1]), 
        .QN(N637) );
  DFFRX2TF \gr_reg[4][2]  ( .D(N980), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[2]), 
        .QN(N636) );
  DFFRX2TF \gr_reg[4][0]  ( .D(N982), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[0]), 
        .QN(N638) );
  DFFSX2TF \pc_reg[6]  ( .D(N817), .CK(CLK), .SN(RST_N), .QN(I_ADDR[7]) );
  DFFSX2TF \pc_reg[4]  ( .D(N822), .CK(CLK), .SN(RST_N), .QN(I_ADDR[5]) );
  DFFSX2TF \pc_reg[1]  ( .D(N825), .CK(CLK), .SN(RST_N), .QN(I_ADDR[2]) );
  DFFSX2TF \pc_reg[0]  ( .D(N874), .CK(CLK), .SN(RST_N), .QN(I_ADDR[1]) );
  DFFRX2TF \gr_reg[1][0]  ( .D(N1006), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[0]), 
        .QN(N686) );
  DFFRX2TF \gr_reg[1][1]  ( .D(N1005), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[1]), 
        .QN(N685) );
  DFFRX2TF \gr_reg[2][11]  ( .D(N955), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTA[11]), .QN(N659) );
  DFFRX2TF \gr_reg[2][12]  ( .D(N954), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTA[12]), .QN(N658) );
  DFFRX2TF \gr_reg[2][8]  ( .D(N958), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[8]), 
        .QN(N662) );
  DFFRX2TF \gr_reg[2][10]  ( .D(N956), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTA[10]), .QN(N660) );
  DFFRX2TF \gr_reg[2][9]  ( .D(N957), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[9]), 
        .QN(N661) );
  DFFRX2TF \gr_reg[2][5]  ( .D(N993), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[5]), 
        .QN(N665) );
  DFFRX2TF \gr_reg[2][3]  ( .D(N995), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[3]), 
        .QN(N667) );
  DFFRX2TF \gr_reg[1][2]  ( .D(N1004), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[2]), 
        .QN(N684) );
  DFFRX2TF \gr_reg[1][4]  ( .D(N1002), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[4]), 
        .QN(N682) );
  DFFRX2TF \gr_reg[2][1]  ( .D(N997), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[1]), 
        .QN(N669) );
  DFFRX2TF \gr_reg[2][6]  ( .D(N992), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[6]), 
        .QN(N664) );
  DFFRX2TF \gr_reg[2][2]  ( .D(N996), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[2]), 
        .QN(N668) );
  DFFRX2TF \gr_reg[2][7]  ( .D(N991), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[7]), 
        .QN(N663) );
  DFFRX2TF \gr_reg[2][4]  ( .D(N994), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[4]), 
        .QN(N666) );
  DFFRX2TF \gr_reg[2][0]  ( .D(N998), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[0]), 
        .QN(N670) );
  DFFRX2TF \gr_reg[3][3]  ( .D(N987), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[3]), 
        .QN(N651) );
  CMPR32X2TF \sub_x_283_4/U14  ( .A(N219), .B(REG_A[3]), .C(SUB_X_283_4_N14), 
        .CO(SUB_X_283_4_N13), .S(N503) );
  CMPR32X2TF \sub_x_283_4/U13  ( .A(N220), .B(REG_A[4]), .C(SUB_X_283_4_N13), 
        .CO(SUB_X_283_4_N12), .S(N504) );
  CMPR32X2TF \sub_x_283_4/U10  ( .A(N223), .B(REG_A[7]), .C(SUB_X_283_4_N10), 
        .CO(SUB_X_283_4_N9), .S(N507) );
  CMPR32X2TF \sub_x_283_4/U12  ( .A(N221), .B(REG_A[5]), .C(SUB_X_283_4_N12), 
        .CO(SUB_X_283_4_N11), .S(N505) );
  ADDFHX1TF \sub_x_283_4/U4  ( .A(N229), .B(REG_A[13]), .CI(SUB_X_283_4_N4), 
        .CO(SUB_X_283_4_N3), .S(N513) );
  CMPR32X2TF \sub_x_283_4/U16  ( .A(N21), .B(REG_A[1]), .C(SUB_X_283_4_N16), 
        .CO(SUB_X_283_4_N15), .S(N501) );
  CMPR32X2TF \sub_x_283_4/U15  ( .A(N218), .B(REG_A[2]), .C(SUB_X_283_4_N15), 
        .CO(SUB_X_283_4_N14), .S(N502) );
  CMPR32X2TF \add_x_283_3/U12  ( .A(REG_A[5]), .B(REG_B[5]), .C(
        ADD_X_283_3_N12), .CO(ADD_X_283_3_N11), .S(N471) );
  CMPR32X2TF \add_x_283_3/U11  ( .A(REG_A[6]), .B(REG_B[6]), .C(
        ADD_X_283_3_N11), .CO(ADD_X_283_3_N10), .S(N472) );
  CMPR32X2TF \add_x_283_3/U10  ( .A(REG_A[7]), .B(REG_B[7]), .C(
        ADD_X_283_3_N10), .CO(ADD_X_283_3_N9), .S(N473) );
  CMPR32X2TF \add_x_283_3/U3  ( .A(REG_A[14]), .B(REG_B[14]), .C(
        ADD_X_283_3_N3), .CO(ADD_X_283_3_N2), .S(N480) );
  DFFRX2TF \gr_reg[1][5]  ( .D(N1001), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[5]), 
        .QN(N681) );
  DFFNSRX2TF lowest_bit_reg ( .D(N1016), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        N1620), .QN(N160) );
  DFFNSRXLTF \reg_C_reg[9]  ( .D(N518), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N424) );
  DFFNSRXLTF \reg_C_reg[11]  ( .D(N533), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N418) );
  DFFNSRXLTF \reg_C_reg[8]  ( .D(N5090), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N429) );
  DFFNSRXLTF \reg_C_reg[12]  ( .D(N524), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N423) );
  DFFNSRXLTF \reg_C_reg[10]  ( .D(N527), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N421) );
  DFFNSRXLTF \reg_C_reg[13]  ( .D(N530), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N420) );
  DFFNSRXLTF \reg_C_reg[14]  ( .D(N536), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N417) );
  DFFNSRXLTF \reg_C_reg[15]  ( .D(N542), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N412) );
  DFFNSRXLTF is_i_addr_reg ( .D(N114), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        IS_I_ADDR) );
  DFFNSRXLTF dw_reg ( .D(N612), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(D_WE) );
  DFFRX4TF \reg_A_reg[0]  ( .D(N464), .CK(CLK), .RN(RST_N), .Q(REG_A[0]), .QN(
        N243) );
  DFFRX4TF \reg_B_reg[2]  ( .D(N519), .CK(CLK), .RN(RST_N), .Q(REG_B[2]), .QN(
        N218) );
  DFFRX1TF \smdr_reg[5]  ( .D(N484), .CK(CLK), .RN(RST_N), .QN(N615) );
  DFFRX1TF \smdr_reg[13]  ( .D(N4760), .CK(CLK), .RN(RST_N), .QN(N607) );
  DFFRX1TF \smdr_reg[12]  ( .D(N4770), .CK(CLK), .RN(RST_N), .QN(N608) );
  DFFRX1TF \smdr_reg[8]  ( .D(N4810), .CK(CLK), .RN(RST_N), .QN(N6120) );
  DFFRX1TF \smdr_reg[15]  ( .D(N4820), .CK(CLK), .RN(RST_N), .QN(N605) );
  DFFRX1TF \smdr_reg[0]  ( .D(N488), .CK(CLK), .RN(RST_N), .QN(N620) );
  DFFRX1TF \smdr_reg[7]  ( .D(N462), .CK(CLK), .RN(RST_N), .QN(N613) );
  DFFRX1TF \smdr_reg[3]  ( .D(N458), .CK(CLK), .RN(RST_N), .QN(N617) );
  DFFRX1TF \smdr_reg[11]  ( .D(N4780), .CK(CLK), .RN(RST_N), .QN(N609) );
  DFFRX1TF \smdr_reg[1]  ( .D(N487), .CK(CLK), .RN(RST_N), .QN(N619) );
  DFFRX1TF \smdr_reg[6]  ( .D(N483), .CK(CLK), .RN(RST_N), .QN(N614) );
  DFFRX1TF \smdr_reg[4]  ( .D(N485), .CK(CLK), .RN(RST_N), .QN(N616) );
  DFFRX1TF \smdr_reg[14]  ( .D(N4750), .CK(CLK), .RN(RST_N), .QN(N606) );
  DFFRX1TF \smdr_reg[10]  ( .D(N4790), .CK(CLK), .RN(RST_N), .QN(N610) );
  DFFRX1TF \smdr_reg[9]  ( .D(N4800), .CK(CLK), .RN(RST_N), .QN(N611) );
  DFFRX1TF \smdr_reg[2]  ( .D(N486), .CK(CLK), .RN(RST_N), .QN(N618) );
  DFFRX1TF \id_ir_reg[7]  ( .D(N463), .CK(CLK), .RN(RST_N), .QN(N432) );
  DFFRX1TF \id_ir_reg[3]  ( .D(N4700), .CK(CLK), .RN(RST_N), .QN(N431) );
  DFFRX1TF \id_ir_reg[9]  ( .D(N498), .CK(CLK), .RN(RST_N), .Q(N1630), .QN(N22) );
  DFFRX1TF \gr_reg[2][15]  ( .D(N951), .CK(CLK), .RN(RST_N), .QN(N655) );
  DFFRX1TF \gr_reg[2][14]  ( .D(N952), .CK(CLK), .RN(RST_N), .QN(N656) );
  DFFRX1TF \gr_reg[2][13]  ( .D(N953), .CK(CLK), .RN(RST_N), .QN(N657) );
  DFFRX1TF \gr_reg[4][15]  ( .D(N1015), .CK(CLK), .RN(RST_N), .QN(N623) );
  DFFRX1TF \gr_reg[4][14]  ( .D(N936), .CK(CLK), .RN(RST_N), .QN(N624) );
  DFFRX1TF \gr_reg[4][13]  ( .D(N937), .CK(CLK), .RN(RST_N), .QN(N625) );
  DFFRX1TF \gr_reg[4][12]  ( .D(N938), .CK(CLK), .RN(RST_N), .QN(N626) );
  DFFRX1TF \gr_reg[4][11]  ( .D(N939), .CK(CLK), .RN(RST_N), .QN(N627) );
  DFFRX1TF \gr_reg[4][10]  ( .D(N940), .CK(CLK), .RN(RST_N), .QN(N628) );
  DFFRX1TF \gr_reg[1][15]  ( .D(N959), .CK(CLK), .RN(RST_N), .QN(N671) );
  DFFRX1TF \gr_reg[1][14]  ( .D(N960), .CK(CLK), .RN(RST_N), .QN(N672) );
  DFFRX1TF \gr_reg[1][13]  ( .D(N961), .CK(CLK), .RN(RST_N), .QN(N673) );
  DFFRX1TF \gr_reg[1][12]  ( .D(N962), .CK(CLK), .RN(RST_N), .QN(N674) );
  DFFRX1TF \gr_reg[1][11]  ( .D(N963), .CK(CLK), .RN(RST_N), .QN(N675) );
  DFFRX1TF \gr_reg[1][10]  ( .D(N964), .CK(CLK), .RN(RST_N), .QN(N676) );
  DFFRX1TF \gr_reg[1][9]  ( .D(N965), .CK(CLK), .RN(RST_N), .QN(N677) );
  DFFRX1TF \gr_reg[1][8]  ( .D(N966), .CK(CLK), .RN(RST_N), .QN(N678) );
  DFFRX1TF \gr_reg[0][15]  ( .D(N967), .CK(CLK), .RN(RST_N), .QN(N687) );
  DFFRX1TF \gr_reg[0][14]  ( .D(N968), .CK(CLK), .RN(RST_N), .QN(N688) );
  DFFRX1TF \gr_reg[0][13]  ( .D(N969), .CK(CLK), .RN(RST_N), .QN(N689) );
  DFFRX1TF \gr_reg[0][12]  ( .D(N970), .CK(CLK), .RN(RST_N), .QN(N690) );
  DFFRX1TF \gr_reg[0][11]  ( .D(N971), .CK(CLK), .RN(RST_N), .QN(N691) );
  DFFRX1TF \gr_reg[0][10]  ( .D(N972), .CK(CLK), .RN(RST_N), .QN(N692) );
  DFFRX1TF \gr_reg[0][9]  ( .D(N973), .CK(CLK), .RN(RST_N), .QN(N693) );
  DFFRX1TF \gr_reg[0][8]  ( .D(N974), .CK(CLK), .RN(RST_N), .QN(N694) );
  DFFRX1TF \gr_reg[1][7]  ( .D(N999), .CK(CLK), .RN(RST_N), .QN(N679) );
  DFFRX1TF \gr_reg[0][5]  ( .D(N1009), .CK(CLK), .RN(RST_N), .QN(N697) );
  DFFRX1TF \gr_reg[0][0]  ( .D(N1014), .CK(CLK), .RN(RST_N), .QN(N702) );
  DFFRX1TF \gr_reg[0][7]  ( .D(N1007), .CK(CLK), .RN(RST_N), .QN(N695) );
  DFFRX1TF \gr_reg[0][6]  ( .D(N1008), .CK(CLK), .RN(RST_N), .QN(N696) );
  DFFRX1TF \gr_reg[0][4]  ( .D(N1010), .CK(CLK), .RN(RST_N), .QN(N698) );
  DFFRX1TF \gr_reg[0][3]  ( .D(N1011), .CK(CLK), .RN(RST_N), .QN(N699) );
  DFFRX1TF \gr_reg[0][2]  ( .D(N1012), .CK(CLK), .RN(RST_N), .QN(N700) );
  DFFRX1TF \gr_reg[0][1]  ( .D(N1013), .CK(CLK), .RN(RST_N), .QN(N701) );
  DFFSRX2TF \state_reg[2]  ( .D(NEXT_STATE[2]), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(N267), .QN(N564) );
  DFFSRX2TF \reg_A_reg[13]  ( .D(N528), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_A[13]), .QN(N248) );
  DFFSRX2TF \reg_A_reg[11]  ( .D(N531), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_A[11]), .QN(N257) );
  DFFSRX2TF \reg_A_reg[10]  ( .D(N525), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_A[10]), .QN(N251) );
  DFFSRX2TF \reg_A_reg[9]  ( .D(N5160), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_A[9]), .QN(N250) );
  DFFSRX2TF \reg_A_reg[8]  ( .D(N5070), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_A[8]), .QN(N252) );
  DFFSRX2TF \reg_A_reg[7]  ( .D(N461), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_A[7]), .QN(N255) );
  DFFSRX2TF \reg_A_reg[5]  ( .D(N5040), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_A[5]), .QN(N254) );
  DFFSRX2TF \reg_A_reg[2]  ( .D(N4660), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_A[2]), .QN(N256) );
  DFFSRX2TF \state_reg[0]  ( .D(NEXT_STATE[0]), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(STATE[0]), .QN(N244) );
  DFFSRX2TF \reg_A_reg[15]  ( .D(N540), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_A[15]), .QN(N247) );
  DFFSRX2TF \reg_A_reg[14]  ( .D(N534), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_A[14]), .QN(N241) );
  DFFSRX2TF \reg_A_reg[12]  ( .D(N522), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_A[12]), .QN(N253) );
  DFFSRX2TF \reg_A_reg[1]  ( .D(N465), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_A[1]), .QN(N239) );
  DFFSRX2TF \reg_A_reg[3]  ( .D(N457), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_A[3]), .QN(N258) );
  DFFSRX2TF \reg_A_reg[4]  ( .D(N5130), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_A[4]), .QN(N246) );
  DFFSRX2TF \reg_A_reg[6]  ( .D(N5100), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_A[6]), .QN(N249) );
  DFFSRX2TF \reg_B_reg[12]  ( .D(N449), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_B[12]), .QN(N228) );
  DFFSRX2TF \reg_B_reg[15]  ( .D(N443), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_B[15]), .QN(N231) );
  DFFSRX2TF \reg_B_reg[9]  ( .D(N450), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_B[9]), .QN(N225) );
  DFFSRX2TF \reg_B_reg[14]  ( .D(N444), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_B[14]), .QN(N230) );
  DFFSRX2TF \reg_B_reg[11]  ( .D(N445), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_B[11]), .QN(N227) );
  DFFSRX2TF nf_reg ( .D(N442), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(NF), .QN(
        N271) );
  DFFSRX2TF \reg_B_reg[7]  ( .D(N455), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_B[7]), .QN(N223) );
  DFFSRX2TF \reg_B_reg[3]  ( .D(N456), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_B[3]), .QN(N219) );
  DFFSRX2TF \reg_B_reg[6]  ( .D(N452), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_B[6]), .QN(N222) );
  DFFSRX2TF \reg_B_reg[5]  ( .D(N454), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_B[5]), .QN(N221) );
  DFFSRX2TF \reg_B_reg[4]  ( .D(N451), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_B[4]), .QN(N220) );
  DFFSRX2TF \reg_B_reg[10]  ( .D(N447), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_B[10]), .QN(N226) );
  DFFSRX2TF \reg_B_reg[8]  ( .D(N453), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_B[8]), .QN(N224) );
  DFFSRX2TF \reg_B_reg[13]  ( .D(N446), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_B[13]), .QN(N229) );
  DFFSRX2TF zf_reg ( .D(N448), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(ZF), .QN(
        N272) );
  DFFSRX2TF \id_ir_reg[6]  ( .D(N4670), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        N273), .QN(N414) );
  DFFSRX2TF \id_ir_reg[5]  ( .D(N4680), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        N274), .QN(N415) );
  DFFSRX2TF \id_ir_reg[4]  ( .D(N4690), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        N275), .QN(N416) );
  DFFSRX2TF \id_ir_reg[2]  ( .D(N4710), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        OPER3_R3[2]), .QN(N276) );
  DFFSRX2TF \id_ir_reg[0]  ( .D(N4730), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        OPER3_R3[0]), .QN(N265) );
  DFFSRX2TF \id_ir_reg[14]  ( .D(N493), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        CODE_TYPE[3]), .QN(N266) );
  DFFSRX2TF \id_ir_reg[13]  ( .D(N494), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        CODE_TYPE[2]), .QN(N262) );
  DFFSRX2TF \id_ir_reg[12]  ( .D(N495), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        N245), .QN(N23) );
  DFFSRX2TF \id_ir_reg[10]  ( .D(N497), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        \OPER1_R1[2] ), .QN(N264) );
  DFFSRX2TF \id_ir_reg[8]  ( .D(N499), .CK(CLK), .SN(1'b1), .RN(RST_N), .Q(
        N259), .QN(N582) );
  DFFRX1TF \state_reg[1]  ( .D(NEXT_STATE[1]), .CK(CLK), .RN(RST_N), .Q(
        STATE[1]) );
  DFFRX1TF cf_reg ( .D(N4740), .CK(CLK), .RN(RST_N), .Q(CF) );
  DFFRX2TF \gr_reg[1][6]  ( .D(N1000), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[6]), 
        .QN(N680) );
  DFFNSRX2TF \reg_C_reg[5]  ( .D(N5060), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[6]) );
  DFFNSRX2TF \reg_C_reg[3]  ( .D(N460), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[4]) );
  DFFNSRX2TF \reg_C_reg[0]  ( .D(N545), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[1]) );
  DFFNSRX2TF \reg_C_reg[7]  ( .D(N5030), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[8]) );
  DFFNSRX2TF \reg_C_reg[2]  ( .D(N521), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[3]) );
  DFFNSRX2TF \reg_C_reg[6]  ( .D(N5120), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[7]) );
  DFFNSRX2TF \reg_C_reg[4]  ( .D(N5150), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[5]) );
  DFFNSRX2TF \reg_C_reg[1]  ( .D(N539), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[2]) );
  DFFRX2TF \reg_B_reg[1]  ( .D(N537), .CK(CLK), .RN(RST_N), .Q(REG_B[1]), .QN(
        N21) );
  OR3X1TF U3 ( .A(N23), .B(N904), .C(N398), .Y(N839) );
  ADDHXLTF U4 ( .A(REG_B[0]), .B(REG_A[0]), .CO(ADD_X_283_3_N16), .S(N466) );
  NAND2BX1TF U5 ( .AN(REG_A[0]), .B(REG_B[0]), .Y(SUB_X_283_4_N16) );
  INVX2TF U6 ( .A(N726), .Y(N789) );
  NAND3X1TF U7 ( .A(N23), .B(N935), .C(N903), .Y(N829) );
  ADDFHX2TF U8 ( .A(REG_A[11]), .B(REG_B[11]), .CI(ADD_X_283_3_N6), .CO(
        ADD_X_283_3_N5), .S(N477) );
  NAND2X1TF U9 ( .A(N1205), .B(N1204), .Y(N1203) );
  NAND2X1TF U10 ( .A(N562), .B(N244), .Y(N382) );
  OAI22X1TF U11 ( .A0(N1208), .A1(N1185), .B0(N1184), .B1(N1183), .Y(N1186) );
  AOI211X2TF U12 ( .A0(N846), .A1(N759), .B0(N523), .C0(N520), .Y(N1209) );
  ADDFX2TF U13 ( .A(REG_A[15]), .B(REG_B[15]), .CI(ADD_X_283_3_N2), .CO(N482), 
        .S(N481) );
  AOI22X1TF U14 ( .A0(N1188), .A1(D_ADDR[1]), .B0(N175), .B1(IO_DATAINB[0]), 
        .Y(N1) );
  AOI22X1TF U15 ( .A0(N1201), .A1(IO_STATUS[0]), .B0(IO_DATAINA[0]), .B1(N206), 
        .Y(N2) );
  NAND3X1TF U16 ( .A(N1), .B(N1216), .C(N2), .Y(N545) );
  AOI211X1TF U17 ( .A0(REG_A[10]), .A1(N211), .B0(N740), .C0(N705), .Y(N3) );
  NAND2X1TF U18 ( .A(N572), .B(N3), .Y(N535) );
  OA21XLTF U19 ( .A0(I_ADDR[1]), .A1(I_ADDR[2]), .B0(N354), .Y(N4) );
  AOI222XLTF U20 ( .A0(I_ADDR[2]), .A1(N368), .B0(D_ADDR[2]), .B1(N367), .C0(
        N365), .C1(N4), .Y(N825) );
  AOI21X1TF U21 ( .A0(N192), .A1(REG_A[4]), .B0(N739), .Y(N5) );
  NAND3X1TF U22 ( .A(N571), .B(N781), .C(N5), .Y(N759) );
  OA22X1TF U23 ( .A0(N371), .A1(N370), .B0(N380), .B1(N373), .Y(N6) );
  NAND2X1TF U24 ( .A(N1029), .B(START), .Y(N7) );
  OA22X1TF U25 ( .A0(N377), .A1(N374), .B0(STATE[1]), .B1(N7), .Y(N8) );
  NAND4X1TF U26 ( .A(N1188), .B(N381), .C(N6), .D(N8), .Y(NEXT_STATE[0]) );
  OA21XLTF U27 ( .A0(N358), .A1(I_ADDR[5]), .B0(N361), .Y(N9) );
  AOI222XLTF U28 ( .A0(I_ADDR[5]), .A1(N368), .B0(D_ADDR[5]), .B1(N367), .C0(
        N365), .C1(N9), .Y(N822) );
  NOR4XLTF U29 ( .A(N1212), .B(N1203), .C(N1207), .D(N1109), .Y(N10) );
  NOR4XLTF U30 ( .A(N1123), .B(N1103), .C(N1097), .D(N1116), .Y(N11) );
  NOR3X1TF U31 ( .A(N1131), .B(N1160), .C(N1130), .Y(N12) );
  NAND4X1TF U32 ( .A(N10), .B(N11), .C(N12), .D(N1138), .Y(N13) );
  NAND4BX1TF U33 ( .AN(N1041), .B(N1173), .C(N1209), .D(N1184), .Y(N14) );
  OAI2BB2XLTF U34 ( .B0(N13), .B1(N14), .A0N(N1041), .A1N(ZF), .Y(N448) );
  OA21XLTF U35 ( .A0(N366), .A1(I_ADDR[7]), .B0(N364), .Y(N15) );
  AOI222XLTF U36 ( .A0(I_ADDR[7]), .A1(N368), .B0(D_ADDR[7]), .B1(N367), .C0(
        N365), .C1(N15), .Y(N817) );
  AOI21X1TF U37 ( .A0(N192), .A1(REG_A[11]), .B0(N550), .Y(N16) );
  NAND3X1TF U38 ( .A(N549), .B(N596), .C(N16), .Y(N771) );
  OAI22X1TF U39 ( .A0(N1184), .A1(N1185), .B0(N1205), .B1(N1183), .Y(N17) );
  AOI21X1TF U40 ( .A0(IO_DATAINA[14]), .A1(N206), .B0(N17), .Y(N18) );
  OAI21X1TF U41 ( .A0(N170), .A1(N417), .B0(N18), .Y(N536) );
  AOI21X1TF U42 ( .A0(N354), .A1(N280), .B0(N360), .Y(N19) );
  AOI222XLTF U43 ( .A0(I_ADDR[3]), .A1(N368), .B0(N19), .B1(N355), .C0(N367), 
        .C1(D_ADDR[3]), .Y(N824) );
  ADDFHX2TF U44 ( .A(REG_A[12]), .B(REG_B[12]), .CI(ADD_X_283_3_N5), .CO(
        ADD_X_283_3_N4), .S(N478) );
  ADDFHX4TF U45 ( .A(REG_A[9]), .B(REG_B[9]), .CI(ADD_X_283_3_N8), .CO(
        ADD_X_283_3_N7), .S(N475) );
  AOI22X4TF U46 ( .A0(N1215), .A1(N1214), .B0(N1213), .B1(N1212), .Y(N1216) );
  INVXLTF U47 ( .A(N23), .Y(N24) );
  AOI22XLTF U48 ( .A0(N315), .A1(N328), .B0(N680), .B1(N314), .Y(N1000) );
  NAND2XLTF U110 ( .A(N192), .B(REG_A[3]), .Y(N556) );
  NAND2XLTF U111 ( .A(N211), .B(REG_A[11]), .Y(N392) );
  NAND2XLTF U112 ( .A(N726), .B(N219), .Y(N5050) );
  OR3X1TF U113 ( .A(REG_B[2]), .B(REG_B[3]), .C(N829), .Y(N853) );
  AO22X1TF U114 ( .A0(\OPER1_R1[2] ), .A1(N914), .B0(N913), .B1(N273), .Y(
        N1178) );
  OR3X1TF U115 ( .A(N178), .B(N934), .C(N933), .Y(N1200) );
  AO22X1TF U116 ( .A0(N928), .A1(N914), .B0(N416), .B1(N911), .Y(N1176) );
  INVX2TF U117 ( .A(N837), .Y(N186) );
  NAND2XLTF U118 ( .A(N192), .B(REG_A[2]), .Y(N780) );
  NAND3XLTF U119 ( .A(N373), .B(N381), .C(N372), .Y(NEXT_STATE[1]) );
  OR4X2TF U120 ( .A(N23), .B(N924), .C(N923), .D(N922), .Y(N1084) );
  INVX2TF U121 ( .A(N593), .Y(N158) );
  NAND2XLTF U122 ( .A(N593), .B(REG_A[6]), .Y(N594) );
  NAND3X2TF U123 ( .A(STATE[0]), .B(N405), .C(N263), .Y(N310) );
  CLKINVX1TF U124 ( .A(N904), .Y(N385) );
  OR2X2TF U125 ( .A(REG_B[0]), .B(N21), .Y(N793) );
  OR3X2TF U126 ( .A(N564), .B(STATE[1]), .C(N382), .Y(N1188) );
  OAI31X2TF U127 ( .A0(REG_B[3]), .A1(N789), .A2(N756), .B0(N532), .Y(N546) );
  AOI21X2TF U128 ( .A0(N479), .A1(N187), .B0(N800), .Y(N802) );
  OAI21X1TF U129 ( .A0(N634), .A1(N214), .B0(N1076), .Y(N485) );
  OAI21X1TF U130 ( .A0(N637), .A1(N210), .B0(N1169), .Y(N537) );
  OAI21X1TF U131 ( .A0(N633), .A1(N213), .B0(N1073), .Y(N484) );
  OAI21X1TF U132 ( .A0(N636), .A1(N210), .B0(N1137), .Y(N519) );
  OAI21XLTF U133 ( .A0(N680), .A1(N1182), .B0(N1115), .Y(N5100) );
  OAI21X1TF U134 ( .A0(N638), .A1(N210), .B0(N1198), .Y(N543) );
  OAI21X1TF U135 ( .A0(N632), .A1(N214), .B0(N1070), .Y(N483) );
  OAI21X1TF U136 ( .A0(N623), .A1(N214), .B0(N1067), .Y(N4820) );
  OAI21X1TF U137 ( .A0(N630), .A1(N213), .B0(N1064), .Y(N4810) );
  OAI21X1TF U138 ( .A0(N629), .A1(N214), .B0(N1061), .Y(N4800) );
  OAI21X1TF U139 ( .A0(N628), .A1(N214), .B0(N1058), .Y(N4790) );
  OAI21X1TF U140 ( .A0(N627), .A1(N214), .B0(N1055), .Y(N4780) );
  OAI21X1TF U141 ( .A0(N624), .A1(N214), .B0(N1046), .Y(N4750) );
  OAI21X1TF U142 ( .A0(N626), .A1(N213), .B0(N1052), .Y(N4770) );
  OAI21X1TF U143 ( .A0(N625), .A1(N213), .B0(N1049), .Y(N4760) );
  OAI21X1TF U144 ( .A0(N636), .A1(N214), .B0(N1079), .Y(N486) );
  OAI21X1TF U145 ( .A0(N638), .A1(N214), .B0(N1090), .Y(N488) );
  OAI21X1TF U146 ( .A0(N637), .A1(N214), .B0(N1082), .Y(N487) );
  OAI21X1TF U147 ( .A0(N635), .A1(N210), .B0(N895), .Y(N456) );
  AOI211X1TF U148 ( .A0(N1089), .A1(IO_DATAOUTB[5]), .B0(N1072), .C0(N1071), 
        .Y(N1073) );
  AOI211X1TF U149 ( .A0(N204), .A1(IO_DATAOUTB[6]), .B0(N1069), .C0(N1068), 
        .Y(N1070) );
  AOI211X1TF U150 ( .A0(N1089), .A1(IO_DATAOUTB[2]), .B0(N1078), .C0(N1077), 
        .Y(N1079) );
  AOI211X1TF U151 ( .A0(N1089), .A1(N278), .B0(N1045), .C0(N1044), .Y(N1046)
         );
  AOI211X1TF U152 ( .A0(N204), .A1(IO_DATAOUTB[4]), .B0(N1075), .C0(N1074), 
        .Y(N1076) );
  AOI211X1TF U153 ( .A0(N1089), .A1(IO_DATAOUTB[9]), .B0(N1060), .C0(N1059), 
        .Y(N1061) );
  AOI211X1TF U154 ( .A0(N1089), .A1(IO_DATAOUTB[10]), .B0(N1057), .C0(N1056), 
        .Y(N1058) );
  AOI211X1TF U155 ( .A0(N1089), .A1(IO_DATAOUTB[0]), .B0(N1088), .C0(N1087), 
        .Y(N1090) );
  AOI211X1TF U156 ( .A0(N204), .A1(IO_DATAOUTB[11]), .B0(N1054), .C0(N1053), 
        .Y(N1055) );
  AOI211X1TF U157 ( .A0(N1089), .A1(IO_DATAOUTB[8]), .B0(N1063), .C0(N1062), 
        .Y(N1064) );
  AOI211X1TF U158 ( .A0(N204), .A1(IO_DATAOUTB[1]), .B0(N1081), .C0(N1080), 
        .Y(N1082) );
  AOI211X1TF U159 ( .A0(N1089), .A1(N279), .B0(N1066), .C0(N1065), .Y(N1067)
         );
  AOI211X1TF U160 ( .A0(N1089), .A1(IO_DATAOUTB[12]), .B0(N1051), .C0(N1050), 
        .Y(N1052) );
  AOI22X1TF U161 ( .A0(N338), .A1(N348), .B0(N675), .B1(N337), .Y(N963) );
  AOI22X1TF U162 ( .A0(N320), .A1(N325), .B0(N651), .B1(N319), .Y(N987) );
  OAI22X1TF U163 ( .A0(N702), .A1(N1086), .B0(N670), .B1(N189), .Y(N1087) );
  AOI22X1TF U164 ( .A0(N344), .A1(N349), .B0(N642), .B1(N342), .Y(N946) );
  AOI22X1TF U165 ( .A0(N338), .A1(N347), .B0(N676), .B1(N337), .Y(N964) );
  AOI22X1TF U166 ( .A0(N340), .A1(N348), .B0(N659), .B1(N339), .Y(N955) );
  AOI22X1TF U167 ( .A0(N317), .A1(N322), .B0(N670), .B1(N316), .Y(N998) );
  AOI22X1TF U168 ( .A0(N340), .A1(N352), .B0(N656), .B1(N339), .Y(N952) );
  OAI22X1TF U169 ( .A0(N697), .A1(N1086), .B0(N665), .B1(N189), .Y(N1071) );
  AOI22X1TF U170 ( .A0(N315), .A1(N326), .B0(N682), .B1(N314), .Y(N1002) );
  AOI22X1TF U171 ( .A0(N338), .A1(N345), .B0(N678), .B1(N337), .Y(N966) );
  AOI22X1TF U172 ( .A0(N315), .A1(N323), .B0(N685), .B1(N314), .Y(N1005) );
  AOI22X1TF U173 ( .A0(N340), .A1(N350), .B0(N657), .B1(N339), .Y(N953) );
  AOI22X1TF U174 ( .A0(N344), .A1(N346), .B0(N645), .B1(N342), .Y(N949) );
  AOI22X1TF U175 ( .A0(N344), .A1(N347), .B0(N644), .B1(N342), .Y(N948) );
  OAI22X1TF U176 ( .A0(N689), .A1(N1086), .B0(N657), .B1(N189), .Y(N1047) );
  AOI22X1TF U177 ( .A0(N340), .A1(N345), .B0(N662), .B1(N339), .Y(N958) );
  OAI22X1TF U178 ( .A0(N690), .A1(N1086), .B0(N658), .B1(N189), .Y(N1050) );
  OAI22X1TF U179 ( .A0(N640), .A1(N201), .B0(N672), .B1(N1191), .Y(N430) );
  AOI22X1TF U180 ( .A0(N344), .A1(N345), .B0(N646), .B1(N342), .Y(N950) );
  AOI22X1TF U181 ( .A0(N344), .A1(N343), .B0(N639), .B1(N342), .Y(N943) );
  AOI22X1TF U182 ( .A0(N317), .A1(N328), .B0(N664), .B1(N316), .Y(N992) );
  AOI22X1TF U183 ( .A0(N320), .A1(N326), .B0(N650), .B1(N319), .Y(N986) );
  OAI22X1TF U184 ( .A0(N642), .A1(N201), .B0(N674), .B1(N1191), .Y(N858) );
  AOI22X1TF U185 ( .A0(N320), .A1(N324), .B0(N652), .B1(N319), .Y(N988) );
  AOI22X1TF U186 ( .A0(N320), .A1(N330), .B0(N647), .B1(N319), .Y(N983) );
  AOI22X1TF U187 ( .A0(N317), .A1(N323), .B0(N669), .B1(N316), .Y(N997) );
  AOI22X1TF U188 ( .A0(N320), .A1(N323), .B0(N653), .B1(N319), .Y(N989) );
  OAI22X1TF U189 ( .A0(N694), .A1(N1086), .B0(N662), .B1(N189), .Y(N1062) );
  AOI22X1TF U190 ( .A0(N317), .A1(N327), .B0(N665), .B1(N316), .Y(N993) );
  OAI22X1TF U191 ( .A0(N641), .A1(N201), .B0(N673), .B1(N1191), .Y(N440) );
  AOI22X1TF U192 ( .A0(N317), .A1(N325), .B0(N667), .B1(N316), .Y(N995) );
  OAI22X1TF U193 ( .A0(N687), .A1(N1086), .B0(N655), .B1(N189), .Y(N1065) );
  AOI22X1TF U194 ( .A0(N340), .A1(N343), .B0(N655), .B1(N339), .Y(N951) );
  OAI22X1TF U195 ( .A0(N196), .A1(N6120), .B0(N678), .B1(N1083), .Y(N1063) );
  AOI22X1TF U196 ( .A0(N335), .A1(N345), .B0(N694), .B1(N334), .Y(N974) );
  AOI22X1TF U197 ( .A0(N313), .A1(N323), .B0(N701), .B1(N312), .Y(N1013) );
  AOI22X1TF U198 ( .A0(N335), .A1(N347), .B0(N692), .B1(N334), .Y(N972) );
  OAI22X1TF U199 ( .A0(N196), .A1(N608), .B0(N674), .B1(N1083), .Y(N1051) );
  AOI22X1TF U200 ( .A0(N335), .A1(N348), .B0(N691), .B1(N334), .Y(N971) );
  OAI22X1TF U201 ( .A0(N195), .A1(N607), .B0(N673), .B1(N1083), .Y(N1048) );
  NAND4XLTF U202 ( .A(N395), .B(N292), .C(N389), .D(N778), .Y(N584) );
  OAI22X1TF U203 ( .A0(N196), .A1(N620), .B0(N686), .B1(N1083), .Y(N1088) );
  AOI22X1TF U204 ( .A0(N313), .A1(N328), .B0(N696), .B1(N312), .Y(N1008) );
  OAI22X1TF U205 ( .A0(N195), .A1(N615), .B0(N681), .B1(N1083), .Y(N1072) );
  AOI22X1TF U206 ( .A0(N313), .A1(N326), .B0(N698), .B1(N312), .Y(N1010) );
  OAI22X1TF U207 ( .A0(N195), .A1(N605), .B0(N671), .B1(N1083), .Y(N1066) );
  OAI22X1TF U208 ( .A0(N627), .A1(N1199), .B0(N659), .B1(N1194), .Y(N435) );
  OAI22X1TF U209 ( .A0(N626), .A1(N1199), .B0(N658), .B1(N1194), .Y(N857) );
  OAI22X1TF U210 ( .A0(N623), .A1(N1199), .B0(N655), .B1(N1194), .Y(N422) );
  AND3X2TF U211 ( .A(OPER3_R3[0]), .B(N411), .C(OPER3_R3[1]), .Y(N1192) );
  NAND4X2TF U212 ( .A(N265), .B(N276), .C(N260), .D(N411), .Y(N1190) );
  NAND2BX2TF U213 ( .AN(N926), .B(N194), .Y(N1083) );
  NAND2BX2TF U214 ( .AN(N927), .B(N194), .Y(N1086) );
  OAI211X1TF U215 ( .A0(N922), .A1(N912), .B0(N915), .C0(N916), .Y(N1175) );
  AND2X2TF U216 ( .A(\OPER1_R1[2] ), .B(N195), .Y(N212) );
  AND2X2TF U217 ( .A(N395), .B(N912), .Y(N835) );
  AND2X2TF U218 ( .A(N928), .B(N194), .Y(N1085) );
  BUFX3TF U219 ( .A(N1202), .Y(N206) );
  OAI211X1TF U220 ( .A0(N23), .A1(N394), .B0(N390), .C0(N389), .Y(N837) );
  INVX1TF U221 ( .A(N808), .Y(N810) );
  INVX1TF U222 ( .A(N886), .Y(N887) );
  OAI211XLTF U223 ( .A0(N383), .A1(N382), .B0(N558), .C0(N381), .Y(
        NEXT_STATE[2]) );
  NAND2X2TF U224 ( .A(N169), .B(N932), .Y(N1183) );
  INVX2TF U225 ( .A(N839), .Y(N165) );
  NAND2XLTF U226 ( .A(REG_B[3]), .B(N726), .Y(N568) );
  AOI22X1TF U227 ( .A0(N198), .A1(REG_A[14]), .B0(N710), .B1(REG_A[13]), .Y(
        N554) );
  AOI32X1TF U228 ( .A0(N1091), .A1(N1620), .A2(N244), .B0(N305), .B1(N1620), 
        .Y(N306) );
  INVX2TF U229 ( .A(N1188), .Y(N169) );
  NAND2XLTF U230 ( .A(N593), .B(REG_A[4]), .Y(N391) );
  INVX2TF U231 ( .A(N779), .Y(N197) );
  NOR2X1TF U232 ( .A(N1640), .B(N582), .Y(N925) );
  INVX1TF U233 ( .A(N1092), .Y(N288) );
  NAND3XLTF U234 ( .A(N905), .B(N903), .C(N245), .Y(N294) );
  INVX1TF U235 ( .A(N374), .Y(N376) );
  INVX2TF U236 ( .A(N1215), .Y(N159) );
  INVX2TF U237 ( .A(N160), .Y(I_ADDR[0]) );
  INVX2TF U238 ( .A(N1630), .Y(N1640) );
  INVX2TF U239 ( .A(N839), .Y(N166) );
  INVX2TF U240 ( .A(N310), .Y(N167) );
  INVX2TF U241 ( .A(N310), .Y(N168) );
  INVX2TF U242 ( .A(N1188), .Y(N170) );
  INVX2TF U243 ( .A(N853), .Y(N171) );
  INVX2TF U244 ( .A(N853), .Y(N172) );
  INVX2TF U245 ( .A(N245), .Y(N173) );
  INVX2TF U246 ( .A(N1200), .Y(N174) );
  INVX2TF U247 ( .A(N1200), .Y(N175) );
  INVX2TF U248 ( .A(N835), .Y(N176) );
  INVX2TF U249 ( .A(N835), .Y(N177) );
  INVX2TF U250 ( .A(N169), .Y(N178) );
  INVX2TF U251 ( .A(N1178), .Y(N179) );
  INVX2TF U252 ( .A(N1178), .Y(N180) );
  INVX2TF U253 ( .A(N1175), .Y(N181) );
  INVX2TF U254 ( .A(N181), .Y(N182) );
  INVX2TF U255 ( .A(N181), .Y(N183) );
  INVX2TF U256 ( .A(N1176), .Y(N184) );
  INVX2TF U257 ( .A(N1176), .Y(N185) );
  INVX2TF U258 ( .A(N186), .Y(N187) );
  INVX2TF U259 ( .A(N186), .Y(N188) );
  INVX2TF U260 ( .A(N1085), .Y(N189) );
  INVX2TF U261 ( .A(N1085), .Y(N190) );
  INVX2TF U262 ( .A(N793), .Y(N191) );
  INVX2TF U263 ( .A(N793), .Y(N192) );
  INVX2TF U264 ( .A(N1084), .Y(N194) );
  INVX2TF U265 ( .A(N1084), .Y(N195) );
  INVX2TF U266 ( .A(N1084), .Y(N196) );
  NOR3BX1TF U267 ( .AN(N386), .B(CODE_TYPE[3]), .C(N262), .Y(N1018) );
  NAND2X1TF U268 ( .A(N245), .B(N240), .Y(N386) );
  NOR2X2TF U269 ( .A(STATE[1]), .B(N267), .Y(N383) );
  AOI22X2TF U270 ( .A0(D_ADDR[4]), .A1(N168), .B0(N378), .B1(D_DATAIN[3]), .Y(
        N325) );
  OAI21X2TF U271 ( .A0(N908), .A1(N907), .B0(N906), .Y(N915) );
  NOR2X1TF U272 ( .A(CODE_TYPE[4]), .B(N398), .Y(N908) );
  AOI22X2TF U273 ( .A0(D_ADDR[6]), .A1(N167), .B0(N378), .B1(D_DATAIN[5]), .Y(
        N327) );
  AOI22X2TF U274 ( .A0(D_ADDR[1]), .A1(N167), .B0(N378), .B1(D_DATAIN[0]), .Y(
        N322) );
  AOI22X2TF U275 ( .A0(D_ADDR[8]), .A1(N168), .B0(N378), .B1(D_DATAIN[7]), .Y(
        N330) );
  AOI22X2TF U276 ( .A0(D_ADDR[3]), .A1(N168), .B0(N378), .B1(D_DATAIN[2]), .Y(
        N324) );
  AOI22X2TF U277 ( .A0(D_ADDR[7]), .A1(N168), .B0(N378), .B1(D_DATAIN[6]), .Y(
        N328) );
  AOI22X2TF U278 ( .A0(D_ADDR[5]), .A1(N168), .B0(N378), .B1(D_DATAIN[4]), .Y(
        N326) );
  AOI2BB2X2TF U279 ( .B0(D_DATAIN[7]), .B1(N333), .A0N(N412), .A1N(N332), .Y(
        N343) );
  AOI2BB2X2TF U280 ( .B0(D_DATAIN[1]), .B1(N333), .A0N(N424), .A1N(N332), .Y(
        N346) );
  AOI2BB2X2TF U281 ( .B0(D_DATAIN[6]), .B1(N333), .A0N(N417), .A1N(N332), .Y(
        N352) );
  AOI2BB2X2TF U282 ( .B0(D_DATAIN[4]), .B1(N333), .A0N(N423), .A1N(N332), .Y(
        N349) );
  AOI2BB2X2TF U283 ( .B0(D_DATAIN[5]), .B1(N333), .A0N(N420), .A1N(N332), .Y(
        N350) );
  AOI2BB2X2TF U284 ( .B0(D_DATAIN[2]), .B1(N333), .A0N(N421), .A1N(N332), .Y(
        N347) );
  AOI2BB2X2TF U285 ( .B0(D_DATAIN[3]), .B1(N333), .A0N(N418), .A1N(N332), .Y(
        N348) );
  NOR3X4TF U286 ( .A(N22), .B(N582), .C(N318), .Y(N320) );
  NOR3X4TF U287 ( .A(N1640), .B(N582), .C(N341), .Y(N344) );
  NOR3X4TF U288 ( .A(N1640), .B(N259), .C(N341), .Y(N340) );
  INVX2TF U289 ( .A(N197), .Y(N198) );
  INVX2TF U290 ( .A(N1022), .Y(N199) );
  INVX2TF U291 ( .A(N1022), .Y(N200) );
  INVX2TF U292 ( .A(N1192), .Y(N201) );
  INVX2TF U293 ( .A(N1192), .Y(N202) );
  CLKBUFX2TF U294 ( .A(N158), .Y(N282) );
  INVX2TF U295 ( .A(N778), .Y(N203) );
  NOR2X1TF U296 ( .A(N904), .B(N933), .Y(N836) );
  INVX2TF U297 ( .A(N1043), .Y(N204) );
  CLKBUFX2TF U298 ( .A(N1190), .Y(N205) );
  NOR2X2TF U299 ( .A(N245), .B(N1170), .Y(N1202) );
  CLKBUFX2TF U300 ( .A(N1177), .Y(N207) );
  CLKBUFX2TF U301 ( .A(N281), .Y(N208) );
  CLKBUFX2TF U302 ( .A(N838), .Y(N281) );
  INVX2TF U303 ( .A(N1021), .Y(N209) );
  INVX2TF U304 ( .A(N883), .Y(N210) );
  NAND2X1TF U305 ( .A(N411), .B(OPER3_R3[2]), .Y(N1199) );
  NOR2X2TF U306 ( .A(N262), .B(N240), .Y(N935) );
  OAI22XLTF U307 ( .A0(N625), .A1(N210), .B0(N657), .B1(N1194), .Y(N439) );
  OAI22XLTF U308 ( .A0(N629), .A1(N1199), .B0(N661), .B1(N1194), .Y(N861) );
  OAI22XLTF U309 ( .A0(N624), .A1(N1199), .B0(N656), .B1(N1194), .Y(N428) );
  OAI22XLTF U310 ( .A0(N643), .A1(N201), .B0(N675), .B1(N1191), .Y(N436) );
  OAI22XLTF U311 ( .A0(N639), .A1(N201), .B0(N671), .B1(N1191), .Y(N425) );
  OAI22XLTF U312 ( .A0(N645), .A1(N201), .B0(N677), .B1(N1191), .Y(N862) );
  NOR2X2TF U313 ( .A(CODE_TYPE[2]), .B(N579), .Y(N905) );
  INVX2TF U314 ( .A(N736), .Y(N211) );
  AOI22X2TF U315 ( .A0(D_ADDR[2]), .A1(N168), .B0(N378), .B1(D_DATAIN[1]), .Y(
        N323) );
  AOI2BB2X2TF U316 ( .B0(D_DATAIN[0]), .B1(N333), .A0N(N429), .A1N(N332), .Y(
        N345) );
  INVX2TF U317 ( .A(N212), .Y(N213) );
  INVX2TF U318 ( .A(N212), .Y(N214) );
  OAI31X4TF U319 ( .A0(N408), .A1(N385), .A2(N908), .B0(N170), .Y(N1041) );
  AOI21XLTF U320 ( .A0(N1092), .A1(N383), .B0(N369), .Y(N373) );
  NOR2X2TF U321 ( .A(N244), .B(N263), .Y(N1092) );
  OAI32X4TF U322 ( .A0(N922), .A1(N901), .A2(N934), .B0(N900), .B1(N922), .Y(
        N914) );
  CLKBUFX2TF U323 ( .A(N1083), .Y(N215) );
  CLKBUFX2TF U324 ( .A(N1086), .Y(N216) );
  NOR3X4TF U325 ( .A(N22), .B(N259), .C(N318), .Y(N317) );
  CLKBUFX2TF U326 ( .A(N1193), .Y(N217) );
  CMPR32X2TF U327 ( .A(REG_A[1]), .B(REG_B[1]), .C(ADD_X_283_3_N16), .CO(
        ADD_X_283_3_N15), .S(N467) );
  CMPR32X2TF U328 ( .A(REG_A[4]), .B(REG_B[4]), .C(ADD_X_283_3_N13), .CO(
        ADD_X_283_3_N12), .S(N470) );
  CMPR32X2TF U329 ( .A(REG_A[13]), .B(REG_B[13]), .C(ADD_X_283_3_N4), .CO(
        ADD_X_283_3_N3), .S(N479) );
  ADDFHX4TF U330 ( .A(REG_A[10]), .B(REG_B[10]), .CI(ADD_X_283_3_N7), .CO(
        ADD_X_283_3_N6), .S(N476) );
  ADDFHX2TF U331 ( .A(REG_A[3]), .B(REG_B[3]), .CI(ADD_X_283_3_N14), .CO(
        ADD_X_283_3_N13), .S(N469) );
  ADDFHX2TF U332 ( .A(REG_A[2]), .B(REG_B[2]), .CI(ADD_X_283_3_N15), .CO(
        ADD_X_283_3_N14), .S(N468) );
  ADDFHX2TF U333 ( .A(REG_A[8]), .B(REG_B[8]), .CI(ADD_X_283_3_N9), .CO(
        ADD_X_283_3_N8), .S(N474) );
  XOR2X1TF U334 ( .A(REG_A[0]), .B(REG_B[0]), .Y(N500) );
  INVX2TF U335 ( .A(SUB_X_283_4_N1), .Y(N516) );
  CMPR32X2TF U336 ( .A(N228), .B(REG_A[12]), .C(SUB_X_283_4_N5), .CO(
        SUB_X_283_4_N4), .S(N512) );
  CMPR32X2TF U337 ( .A(N222), .B(REG_A[6]), .C(SUB_X_283_4_N11), .CO(
        SUB_X_283_4_N10), .S(N506) );
  ADDFHX4TF U338 ( .A(N226), .B(REG_A[10]), .CI(SUB_X_283_4_N7), .CO(
        SUB_X_283_4_N6), .S(N510) );
  ADDFHX4TF U339 ( .A(N227), .B(REG_A[11]), .CI(SUB_X_283_4_N6), .CO(
        SUB_X_283_4_N5), .S(N511) );
  ADDFHX4TF U340 ( .A(N231), .B(REG_A[15]), .CI(SUB_X_283_4_N2), .CO(
        SUB_X_283_4_N1), .S(N515) );
  ADDFHX2TF U341 ( .A(N230), .B(REG_A[14]), .CI(SUB_X_283_4_N3), .CO(
        SUB_X_283_4_N2), .S(N514) );
  ADDFHX4TF U342 ( .A(N224), .B(REG_A[8]), .CI(SUB_X_283_4_N9), .CO(
        SUB_X_283_4_N8), .S(N508) );
  ADDFHX4TF U343 ( .A(N225), .B(REG_A[9]), .CI(SUB_X_283_4_N8), .CO(
        SUB_X_283_4_N7), .S(N509) );
  AOI22X4TF U344 ( .A0(N514), .A1(N281), .B0(N480), .B1(N187), .Y(N532) );
  XNOR2X4TF U345 ( .A(N1211), .B(N1210), .Y(N1214) );
  AOI22X4TF U346 ( .A0(N1209), .A1(N1208), .B0(N1207), .B1(N1206), .Y(N1210)
         );
  NAND4X6TF U347 ( .A(N404), .B(N403), .C(N402), .D(N401), .Y(N1207) );
  NOR4BX4TF U348 ( .AN(N548), .B(N547), .C(N546), .D(N544), .Y(N1184) );
  AOI22X4TF U349 ( .A0(N515), .A1(N208), .B0(N481), .B1(N188), .Y(N404) );
  OAI22X1TF U350 ( .A0(N1041), .A1(N1208), .B0(N1042), .B1(N271), .Y(N442) );
  NOR3X2TF U351 ( .A(N173), .B(N398), .C(N923), .Y(N726) );
  NOR2X1TF U352 ( .A(N262), .B(N386), .Y(N406) );
  NOR2X2TF U353 ( .A(REG_B[1]), .B(N20), .Y(N779) );
  AOI221XLTF U354 ( .A0(CODE_TYPE[4]), .A1(N245), .B0(N934), .B1(N23), .C0(
        N240), .Y(N308) );
  AOI21X1TF U355 ( .A0(STATE[0]), .A1(N405), .B0(N562), .Y(N305) );
  OAI21X1TF U356 ( .A0(N935), .A1(N902), .B0(N903), .Y(N407) );
  AOI32X1TF U357 ( .A0(N935), .A1(N245), .A2(CF), .B0(N23), .B1(N295), .Y(N296) );
  AO21X1TF U358 ( .A0(N1215), .A1(N1212), .B0(N1174), .Y(N539) );
  OAI211X1TF U359 ( .A0(N790), .A1(N789), .B0(N788), .C0(N787), .Y(N1212) );
  CLKINVX4TF U360 ( .A(N1207), .Y(N1208) );
  AOI222XLTF U361 ( .A0(N777), .A1(N827), .B0(N776), .B1(N818), .C0(N807), 
        .C1(N826), .Y(N790) );
  NOR2X2TF U362 ( .A(CODE_TYPE[4]), .B(CODE_TYPE[3]), .Y(N903) );
  AOI31X1TF U363 ( .A0(N383), .A1(START), .A2(N244), .B0(N168), .Y(N290) );
  NAND3BX2TF U364 ( .AN(N409), .B(N1189), .C(N876), .Y(N1193) );
  NAND2X1TF U365 ( .A(N336), .B(N264), .Y(N341) );
  NAND2X1TF U366 ( .A(N264), .B(N321), .Y(N318) );
  NOR2X1TF U367 ( .A(N173), .B(CODE_TYPE[2]), .Y(N902) );
  NOR2X1TF U368 ( .A(CODE_TYPE[3]), .B(N242), .Y(N1017) );
  NAND2X1TF U369 ( .A(N867), .B(N409), .Y(N413) );
  INVX2TF U370 ( .A(N1021), .Y(N1182) );
  AOI21X1TF U371 ( .A0(N309), .A1(N332), .B0(N310), .Y(N336) );
  OAI22X1TF U372 ( .A0(N310), .A1(N332), .B0(N309), .B1(N311), .Y(N321) );
  NAND3X1TF U373 ( .A(N579), .B(N903), .C(N902), .Y(N309) );
  NAND2X1TF U374 ( .A(N405), .B(N1092), .Y(N311) );
  INVX2TF U375 ( .A(N289), .Y(N405) );
  NAND2X1TF U376 ( .A(N267), .B(STATE[1]), .Y(N289) );
  NOR3X4TF U377 ( .A(REG_B[2]), .B(REG_B[3]), .C(N789), .Y(N840) );
  OAI21X1TF U378 ( .A0(N562), .A1(N405), .B0(N290), .Y(N162) );
  INVX2TF U379 ( .A(N1043), .Y(N1089) );
  NAND2X1TF U380 ( .A(N925), .B(N194), .Y(N1043) );
  NOR2BX2TF U381 ( .AN(N336), .B(N927), .Y(N335) );
  NOR2X2TF U382 ( .A(N926), .B(N341), .Y(N338) );
  NOR2BX2TF U383 ( .AN(N321), .B(N927), .Y(N313) );
  NAND3X1TF U384 ( .A(N582), .B(N1640), .C(N264), .Y(N927) );
  NOR2X2TF U385 ( .A(N926), .B(N318), .Y(N315) );
  NAND2X1TF U386 ( .A(N1640), .B(N259), .Y(N926) );
  INVX2TF U387 ( .A(N311), .Y(N378) );
  INVX2TF U388 ( .A(N1213), .Y(N1185) );
  AOI211X4TF U389 ( .A0(REG_A[12]), .A1(N834), .B0(N833), .C0(N832), .Y(N1204)
         );
  AOI211X4TF U390 ( .A0(N513), .A1(N281), .B0(N805), .C0(N804), .Y(N1205) );
  NOR2X1TF U391 ( .A(N242), .B(N266), .Y(N899) );
  NAND3X1TF U392 ( .A(CODE_TYPE[2]), .B(N173), .C(N240), .Y(N933) );
  AO22X1TF U393 ( .A0(N293), .A1(N482), .B0(N516), .B1(N208), .Y(N585) );
  NAND2X1TF U394 ( .A(N267), .B(N1092), .Y(N381) );
  AOI222XLTF U395 ( .A0(N304), .A1(N365), .B0(I_ADDR[8]), .B1(N368), .C0(
        D_ADDR[8]), .C1(N367), .Y(N873) );
  NOR2X1TF U396 ( .A(N364), .B(N270), .Y(N371) );
  NAND2X1TF U397 ( .A(N899), .B(N299), .Y(N302) );
  NAND2X1TF U398 ( .A(N366), .B(I_ADDR[7]), .Y(N364) );
  INVX2TF U399 ( .A(N1096), .Y(N1095) );
  NAND2X2TF U400 ( .A(N1092), .B(N1091), .Y(N1096) );
  INVX2TF U401 ( .A(N1040), .Y(N1039) );
  NAND2X2TF U402 ( .A(N1029), .B(N1091), .Y(N1040) );
  INVX2TF U403 ( .A(N382), .Y(N1029) );
  INVX2TF U404 ( .A(N340), .Y(N339) );
  INVX2TF U405 ( .A(N335), .Y(N334) );
  INVX2TF U406 ( .A(N338), .Y(N337) );
  INVX2TF U407 ( .A(N344), .Y(N342) );
  INVX2TF U408 ( .A(N309), .Y(N333) );
  INVX2TF U409 ( .A(N351), .Y(N353) );
  INVX2TF U410 ( .A(N317), .Y(N316) );
  INVX2TF U411 ( .A(N313), .Y(N312) );
  INVX2TF U412 ( .A(N320), .Y(N319) );
  INVX2TF U413 ( .A(N315), .Y(N314) );
  INVX2TF U414 ( .A(N329), .Y(N331) );
  AND2X2TF U415 ( .A(STATE[1]), .B(N564), .Y(N1091) );
  NAND2X1TF U416 ( .A(N383), .B(N1092), .Y(N377) );
  NAND2X1TF U417 ( .A(N211), .B(REG_A[15]), .Y(N849) );
  NAND2X1TF U418 ( .A(N211), .B(REG_A[5]), .Y(N553) );
  INVX2TF U419 ( .A(N836), .Y(N778) );
  NAND2X1TF U420 ( .A(N191), .B(REG_A[5]), .Y(N721) );
  NAND2X1TF U421 ( .A(N191), .B(REG_A[8]), .Y(N572) );
  AOI21X1TF U422 ( .A0(N710), .A1(REG_A[2]), .B0(N5010), .Y(N567) );
  NAND2X1TF U423 ( .A(N710), .B(REG_A[6]), .Y(N571) );
  NAND2X1TF U424 ( .A(N710), .B(REG_A[0]), .Y(N816) );
  AOI211X1TF U425 ( .A0(CODE_TYPE[2]), .A1(N386), .B0(CODE_TYPE[3]), .C0(N896), 
        .Y(N388) );
  AOI211X1TF U426 ( .A0(N1017), .A1(N406), .B0(N932), .C0(N165), .Y(N395) );
  NOR2X1TF U427 ( .A(N923), .B(N933), .Y(N932) );
  NOR2X1TF U428 ( .A(N286), .B(N208), .Y(N292) );
  AOI21X1TF U429 ( .A0(N380), .A1(N379), .B0(N378), .Y(N558) );
  OAI21X1TF U430 ( .A0(N377), .A1(N376), .B0(N375), .Y(N379) );
  OAI31X1TF U431 ( .A0(N245), .A1(N924), .A2(N923), .B0(N167), .Y(N370) );
  NOR2X1TF U432 ( .A(IO_STATUS[0]), .B(IO_STATUS[1]), .Y(N380) );
  OAI21X1TF U433 ( .A0(N651), .A1(N1043), .B0(N931), .Y(N458) );
  AOI211X1TF U434 ( .A0(N212), .A1(IO_OFFSET[3]), .B0(N930), .C0(N929), .Y(
        N931) );
  OAI22X1TF U435 ( .A0(N699), .A1(N216), .B0(N667), .B1(N190), .Y(N929) );
  OAI22X1TF U436 ( .A0(N196), .A1(N617), .B0(N683), .B1(N215), .Y(N930) );
  OAI21X1TF U437 ( .A0(N647), .A1(N1043), .B0(N1028), .Y(N462) );
  AOI211X1TF U438 ( .A0(N212), .A1(IO_OFFSET[7]), .B0(N1027), .C0(N1026), .Y(
        N1028) );
  OAI22X1TF U439 ( .A0(N695), .A1(N216), .B0(N663), .B1(N190), .Y(N1026) );
  OAI22X1TF U440 ( .A0(N195), .A1(N613), .B0(N679), .B1(N215), .Y(N1027) );
  AOI211X1TF U441 ( .A0(N1089), .A1(N277), .B0(N1048), .C0(N1047), .Y(N1049)
         );
  OAI22X1TF U442 ( .A0(N692), .A1(N216), .B0(N660), .B1(N189), .Y(N1056) );
  OAI22X1TF U443 ( .A0(N196), .A1(N610), .B0(N676), .B1(N215), .Y(N1057) );
  OAI22X1TF U444 ( .A0(N688), .A1(N216), .B0(N656), .B1(N189), .Y(N1044) );
  OAI22X1TF U445 ( .A0(N195), .A1(N606), .B0(N672), .B1(N215), .Y(N1045) );
  OAI22X1TF U446 ( .A0(N693), .A1(N216), .B0(N661), .B1(N190), .Y(N1059) );
  OAI22X1TF U447 ( .A0(N196), .A1(N611), .B0(N677), .B1(N215), .Y(N1060) );
  OAI22X1TF U448 ( .A0(N700), .A1(N216), .B0(N668), .B1(N190), .Y(N1077) );
  OAI22X1TF U449 ( .A0(N195), .A1(N618), .B0(N684), .B1(N215), .Y(N1078) );
  OAI22X1TF U450 ( .A0(N691), .A1(N216), .B0(N659), .B1(N190), .Y(N1053) );
  OAI22X1TF U451 ( .A0(N195), .A1(N609), .B0(N675), .B1(N215), .Y(N1054) );
  OAI22X1TF U452 ( .A0(N701), .A1(N216), .B0(N669), .B1(N190), .Y(N1080) );
  OAI22X1TF U453 ( .A0(N196), .A1(N619), .B0(N685), .B1(N215), .Y(N1081) );
  OAI22X1TF U454 ( .A0(N696), .A1(N216), .B0(N664), .B1(N190), .Y(N1068) );
  OAI22X1TF U455 ( .A0(N196), .A1(N614), .B0(N680), .B1(N215), .Y(N1069) );
  OAI22X1TF U456 ( .A0(N698), .A1(N216), .B0(N666), .B1(N190), .Y(N1074) );
  OAI22X1TF U457 ( .A0(N195), .A1(N616), .B0(N682), .B1(N215), .Y(N1075) );
  INVX2TF U458 ( .A(N1041), .Y(N1042) );
  OAI21X1TF U459 ( .A0(N631), .A1(N210), .B0(N891), .Y(N455) );
  NOR3X1TF U460 ( .A(N890), .B(N889), .C(N888), .Y(N891) );
  OAI22X1TF U461 ( .A0(N663), .A1(N284), .B0(N223), .B1(N1193), .Y(N888) );
  OAI22X1TF U462 ( .A0(N647), .A1(N202), .B0(N679), .B1(N283), .Y(N889) );
  OAI22X1TF U463 ( .A0(N432), .A1(N887), .B0(N695), .B1(N1190), .Y(N890) );
  NOR3X1TF U464 ( .A(N894), .B(N893), .C(N892), .Y(N895) );
  OAI22X1TF U465 ( .A0(N667), .A1(N284), .B0(N219), .B1(N1193), .Y(N892) );
  OAI22X1TF U466 ( .A0(N651), .A1(N201), .B0(N683), .B1(N283), .Y(N893) );
  OAI22X1TF U467 ( .A0(N699), .A1(N205), .B0(N431), .B1(N1189), .Y(N894) );
  OAI21X1TF U468 ( .A0(N230), .A1(N1193), .B0(N434), .Y(N444) );
  NOR3X1TF U469 ( .A(N433), .B(N430), .C(N428), .Y(N434) );
  OAI22X1TF U470 ( .A0(N688), .A1(N1190), .B0(N414), .B1(N876), .Y(N433) );
  OAI21X1TF U471 ( .A0(N225), .A1(N217), .B0(N864), .Y(N450) );
  NOR3X1TF U472 ( .A(N863), .B(N862), .C(N861), .Y(N864) );
  OAI22X1TF U473 ( .A0(N693), .A1(N1190), .B0(N260), .B1(N876), .Y(N863) );
  OAI21X1TF U474 ( .A0(N228), .A1(N217), .B0(N860), .Y(N449) );
  NOR3X1TF U475 ( .A(N859), .B(N858), .C(N857), .Y(N860) );
  OAI22X1TF U476 ( .A0(N690), .A1(N1190), .B0(N416), .B1(N876), .Y(N859) );
  OAI21X1TF U477 ( .A0(N226), .A1(N217), .B0(N5000), .Y(N447) );
  NOR3X1TF U478 ( .A(N491), .B(N490), .C(N489), .Y(N5000) );
  OAI22X1TF U479 ( .A0(N628), .A1(N210), .B0(N660), .B1(N284), .Y(N489) );
  OAI22X1TF U480 ( .A0(N644), .A1(N202), .B0(N676), .B1(N283), .Y(N490) );
  OAI22X1TF U481 ( .A0(N692), .A1(N1190), .B0(N276), .B1(N876), .Y(N491) );
  OAI21X1TF U482 ( .A0(N231), .A1(N217), .B0(N427), .Y(N443) );
  NOR3X1TF U483 ( .A(N426), .B(N425), .C(N422), .Y(N427) );
  OAI22X1TF U484 ( .A0(N687), .A1(N1190), .B0(N432), .B1(N876), .Y(N426) );
  OAI21X1TF U485 ( .A0(N227), .A1(N217), .B0(N438), .Y(N445) );
  NOR3X1TF U486 ( .A(N437), .B(N436), .C(N435), .Y(N438) );
  OAI22X1TF U487 ( .A0(N691), .A1(N205), .B0(N431), .B1(N876), .Y(N437) );
  OAI21X1TF U488 ( .A0(N229), .A1(N217), .B0(N459), .Y(N446) );
  NOR3X1TF U489 ( .A(N441), .B(N440), .C(N439), .Y(N459) );
  OAI22X1TF U490 ( .A0(N689), .A1(N205), .B0(N415), .B1(N876), .Y(N441) );
  OAI21X1TF U491 ( .A0(N224), .A1(N217), .B0(N880), .Y(N453) );
  NOR3X1TF U492 ( .A(N879), .B(N878), .C(N877), .Y(N880) );
  OAI22X1TF U493 ( .A0(N630), .A1(N210), .B0(N662), .B1(N284), .Y(N877) );
  OAI22X1TF U494 ( .A0(N646), .A1(N202), .B0(N678), .B1(N283), .Y(N878) );
  OAI22X1TF U495 ( .A0(N694), .A1(N205), .B0(N265), .B1(N876), .Y(N879) );
  NOR3X1TF U496 ( .A(N1136), .B(N1135), .C(N1134), .Y(N1137) );
  OAI22X1TF U497 ( .A0(N668), .A1(N284), .B0(N218), .B1(N1193), .Y(N1134) );
  OAI22X1TF U498 ( .A0(N652), .A1(N201), .B0(N684), .B1(N283), .Y(N1135) );
  OAI22X1TF U499 ( .A0(N700), .A1(N1190), .B0(N276), .B1(N1189), .Y(N1136) );
  NOR3X1TF U500 ( .A(N1197), .B(N1196), .C(N1195), .Y(N1198) );
  OAI22X1TF U501 ( .A0(N670), .A1(N284), .B0(N20), .B1(N1193), .Y(N1195) );
  OAI22X1TF U502 ( .A0(N654), .A1(N202), .B0(N686), .B1(N283), .Y(N1196) );
  OAI22X1TF U503 ( .A0(N702), .A1(N1190), .B0(N265), .B1(N1189), .Y(N1197) );
  NOR3X1TF U504 ( .A(N1168), .B(N1167), .C(N1166), .Y(N1169) );
  OAI22X1TF U505 ( .A0(N669), .A1(N284), .B0(N21), .B1(N1193), .Y(N1166) );
  OAI22X1TF U506 ( .A0(N653), .A1(N202), .B0(N685), .B1(N283), .Y(N1167) );
  OAI22X1TF U507 ( .A0(N701), .A1(N1190), .B0(N260), .B1(N1189), .Y(N1168) );
  OAI211X1TF U508 ( .A0(N698), .A1(N205), .B0(N869), .C0(N868), .Y(N451) );
  AOI211X1TF U509 ( .A0(N883), .A1(IO_OFFSET[4]), .B0(N866), .C0(N865), .Y(
        N869) );
  OAI22X1TF U510 ( .A0(N666), .A1(N284), .B0(N220), .B1(N1193), .Y(N865) );
  OAI22X1TF U511 ( .A0(N650), .A1(N202), .B0(N682), .B1(N283), .Y(N866) );
  OAI211X1TF U512 ( .A0(N697), .A1(N205), .B0(N885), .C0(N884), .Y(N454) );
  AOI211X1TF U513 ( .A0(N883), .A1(IO_OFFSET[5]), .B0(N882), .C0(N881), .Y(
        N885) );
  OAI22X1TF U514 ( .A0(N665), .A1(N284), .B0(N221), .B1(N1193), .Y(N881) );
  OAI22X1TF U515 ( .A0(N649), .A1(N202), .B0(N681), .B1(N283), .Y(N882) );
  OAI211X1TF U516 ( .A0(N696), .A1(N205), .B0(N875), .C0(N872), .Y(N452) );
  NOR2X1TF U517 ( .A(N867), .B(N922), .Y(N886) );
  AOI211X1TF U518 ( .A0(N883), .A1(IO_OFFSET[6]), .B0(N871), .C0(N870), .Y(
        N875) );
  OAI22X1TF U519 ( .A0(N664), .A1(N284), .B0(N222), .B1(N1193), .Y(N870) );
  NAND2X2TF U520 ( .A(N408), .B(N906), .Y(N876) );
  NOR2X1TF U521 ( .A(OPER3_R3[0]), .B(N413), .Y(N419) );
  OAI22X1TF U522 ( .A0(N648), .A1(N202), .B0(N680), .B1(N283), .Y(N871) );
  NOR2X1TF U523 ( .A(OPER3_R3[1]), .B(N413), .Y(N410) );
  INVX2TF U524 ( .A(N1199), .Y(N883) );
  INVX2TF U525 ( .A(N413), .Y(N411) );
  AOI211X1TF U526 ( .A0(N266), .A1(N933), .B0(N922), .C0(CODE_TYPE[4]), .Y(
        N409) );
  AOI211X1TF U527 ( .A0(CODE_TYPE[4]), .A1(N406), .B0(N899), .C0(N897), .Y(
        N867) );
  OAI21X1TF U528 ( .A0(N651), .A1(N1022), .B0(N921), .Y(N457) );
  AOI211X1TF U529 ( .A0(IO_CONTROL[3]), .A1(N1021), .B0(N920), .C0(N919), .Y(
        N921) );
  OAI21X1TF U530 ( .A0(N675), .A1(N1182), .B0(N1159), .Y(N531) );
  AOI211X1TF U531 ( .A0(IO_DATAOUTB[11]), .A1(N199), .B0(N1158), .C0(N1157), 
        .Y(N1159) );
  OAI21X1TF U532 ( .A0(N677), .A1(N1182), .B0(N1129), .Y(N5160) );
  AOI211X1TF U533 ( .A0(IO_DATAOUTB[9]), .A1(N199), .B0(N1128), .C0(N1127), 
        .Y(N1129) );
  OAI21X1TF U534 ( .A0(N684), .A1(N1182), .B0(N1038), .Y(N4660) );
  AOI211X1TF U535 ( .A0(IO_DATAOUTB[2]), .A1(N199), .B0(N1037), .C0(N1036), 
        .Y(N1038) );
  OAI21X1TF U536 ( .A0(N679), .A1(N1182), .B0(N1025), .Y(N461) );
  AOI211X1TF U537 ( .A0(IO_DATAOUTB[7]), .A1(N199), .B0(N1024), .C0(N1023), 
        .Y(N1025) );
  OAI21X1TF U538 ( .A0(N681), .A1(N1182), .B0(N1102), .Y(N5040) );
  AOI211X1TF U539 ( .A0(IO_DATAOUTB[5]), .A1(N199), .B0(N1101), .C0(N1100), 
        .Y(N1102) );
  OAI21X1TF U540 ( .A0(N676), .A1(N1182), .B0(N1148), .Y(N525) );
  AOI211X1TF U541 ( .A0(IO_DATAOUTB[10]), .A1(N199), .B0(N1147), .C0(N1146), 
        .Y(N1148) );
  OAI21X1TF U542 ( .A0(N673), .A1(N1182), .B0(N1154), .Y(N528) );
  AOI211X1TF U543 ( .A0(N277), .A1(N199), .B0(N1153), .C0(N1152), .Y(N1154) );
  OAI21X1TF U544 ( .A0(N678), .A1(N1182), .B0(N1108), .Y(N5070) );
  AOI211X1TF U545 ( .A0(IO_DATAOUTB[8]), .A1(N199), .B0(N1107), .C0(N1106), 
        .Y(N1108) );
  OAI21X1TF U546 ( .A0(N672), .A1(N1182), .B0(N1165), .Y(N534) );
  AOI211X1TF U547 ( .A0(N278), .A1(N200), .B0(N1164), .C0(N1163), .Y(N1165) );
  AOI211X1TF U548 ( .A0(IO_DATAOUTB[6]), .A1(N200), .B0(N1114), .C0(N1113), 
        .Y(N1115) );
  OAI21X1TF U549 ( .A0(N682), .A1(N209), .B0(N1122), .Y(N5130) );
  AOI211X1TF U550 ( .A0(IO_DATAOUTB[4]), .A1(N200), .B0(N1121), .C0(N1120), 
        .Y(N1122) );
  OAI21X1TF U551 ( .A0(N685), .A1(N209), .B0(N1035), .Y(N465) );
  AOI211X1TF U552 ( .A0(IO_DATAOUTB[1]), .A1(N200), .B0(N1034), .C0(N1033), 
        .Y(N1035) );
  OAI21X1TF U553 ( .A0(N671), .A1(N209), .B0(N1181), .Y(N540) );
  AOI211X1TF U554 ( .A0(N279), .A1(N200), .B0(N1180), .C0(N1179), .Y(N1181) );
  OAI21X1TF U555 ( .A0(N674), .A1(N209), .B0(N1143), .Y(N522) );
  AOI211X1TF U556 ( .A0(IO_DATAOUTB[12]), .A1(N200), .B0(N1142), .C0(N1141), 
        .Y(N1143) );
  OAI21X1TF U557 ( .A0(N686), .A1(N209), .B0(N1032), .Y(N464) );
  AOI211X1TF U558 ( .A0(IO_DATAOUTB[0]), .A1(N200), .B0(N1031), .C0(N1030), 
        .Y(N1032) );
  AOI31X4TF U559 ( .A0(N918), .A1(N415), .A2(N414), .B0(N917), .Y(N1177) );
  NOR2X1TF U560 ( .A(N916), .B(N927), .Y(N917) );
  NOR2X1TF U561 ( .A(N915), .B(N275), .Y(N918) );
  NOR2X1TF U562 ( .A(N415), .B(N915), .Y(N911) );
  NOR2X1TF U563 ( .A(N1640), .B(N259), .Y(N928) );
  AOI22X1TF U564 ( .A0(N925), .A1(N914), .B0(N909), .B1(N274), .Y(N1022) );
  NOR2X1TF U565 ( .A(N416), .B(N915), .Y(N909) );
  INVX2TF U566 ( .A(N914), .Y(N916) );
  AOI211X1TF U567 ( .A0(N899), .A1(N898), .B0(N897), .C0(N896), .Y(N900) );
  NOR2X1TF U568 ( .A(N266), .B(N924), .Y(N897) );
  INVX2TF U569 ( .A(N905), .Y(N924) );
  INVX2TF U570 ( .A(N915), .Y(N913) );
  INVX2TF U571 ( .A(N922), .Y(N906) );
  NAND2X2TF U572 ( .A(N1029), .B(N405), .Y(N922) );
  AOI21X1TF U573 ( .A0(N384), .A1(N901), .B0(N934), .Y(N408) );
  AOI21X1TF U574 ( .A0(D_ADDR[1]), .A1(N367), .B0(N303), .Y(N874) );
  AOI211X1TF U575 ( .A0(N367), .A1(D_ADDR[6]), .B0(N363), .C0(N362), .Y(N821)
         );
  AOI211X1TF U576 ( .A0(N361), .A1(N269), .B0(N366), .C0(N360), .Y(N362) );
  NOR2X1TF U577 ( .A(N269), .B(N359), .Y(N363) );
  AOI211X1TF U578 ( .A0(N367), .A1(D_ADDR[4]), .B0(N357), .C0(N356), .Y(N823)
         );
  AOI211X1TF U579 ( .A0(N355), .A1(N268), .B0(N358), .C0(N360), .Y(N356) );
  NOR2X1TF U580 ( .A(N268), .B(N359), .Y(N357) );
  INVX2TF U581 ( .A(N359), .Y(N368) );
  OAI211X1TF U582 ( .A0(N371), .A1(N310), .B0(N301), .C0(N300), .Y(N359) );
  INVX2TF U583 ( .A(N367), .Y(N300) );
  NOR2X2TF U584 ( .A(N310), .B(N302), .Y(N367) );
  INVX2TF U585 ( .A(N360), .Y(N365) );
  OAI211X1TF U586 ( .A0(CF), .A1(N298), .B0(N297), .C0(N296), .Y(N299) );
  AOI32X1TF U587 ( .A0(N579), .A1(ZF), .A2(N262), .B0(N905), .B1(N272), .Y(
        N297) );
  NOR2X1TF U588 ( .A(N361), .B(N269), .Y(N366) );
  NOR2X1TF U589 ( .A(N355), .B(N268), .Y(N358) );
  AOI22X1TF U590 ( .A0(I_ADDR[0]), .A1(N605), .B0(N613), .B1(N160), .Y(
        D_DATAOUT[7]) );
  AOI22X1TF U591 ( .A0(N1620), .A1(N606), .B0(N614), .B1(N160), .Y(
        D_DATAOUT[6]) );
  AOI22X1TF U592 ( .A0(N1620), .A1(N607), .B0(N615), .B1(N160), .Y(
        D_DATAOUT[5]) );
  AOI22X1TF U593 ( .A0(N1620), .A1(N608), .B0(N616), .B1(N160), .Y(
        D_DATAOUT[4]) );
  AOI22X1TF U594 ( .A0(N1620), .A1(N609), .B0(N617), .B1(N160), .Y(
        D_DATAOUT[3]) );
  AOI22X1TF U595 ( .A0(N1620), .A1(N610), .B0(N618), .B1(N160), .Y(
        D_DATAOUT[2]) );
  AOI22X1TF U596 ( .A0(I_ADDR[0]), .A1(N611), .B0(N619), .B1(N160), .Y(
        D_DATAOUT[1]) );
  AOI22X1TF U597 ( .A0(I_ADDR[0]), .A1(N6120), .B0(N620), .B1(N160), .Y(
        D_DATAOUT[0]) );
  AOI22X1TF U598 ( .A0(N1095), .A1(N1094), .B0(N579), .B1(N1096), .Y(N496) );
  AOI22X1TF U599 ( .A0(N1095), .A1(N1093), .B0(N242), .B1(N1096), .Y(N492) );
  AOI22X1TF U600 ( .A0(N1039), .A1(N1093), .B0(N432), .B1(N1040), .Y(N463) );
  INVX2TF U601 ( .A(I_DATAIN[7]), .Y(N1093) );
  AOI22X1TF U602 ( .A0(N1039), .A1(N1094), .B0(N431), .B1(N1040), .Y(N4700) );
  INVX2TF U603 ( .A(I_DATAIN[3]), .Y(N1094) );
  OAI211X1TF U604 ( .A0(N288), .A1(N267), .B0(N375), .C0(N372), .Y(N114) );
  INVX2TF U605 ( .A(N369), .Y(N375) );
  NOR3X1TF U606 ( .A(STATE[0]), .B(N562), .C(N289), .Y(N369) );
  AOI22X1TF U607 ( .A0(N335), .A1(N352), .B0(N688), .B1(N334), .Y(N968) );
  AOI22X1TF U608 ( .A0(N338), .A1(N346), .B0(N677), .B1(N337), .Y(N965) );
  AOI22X1TF U609 ( .A0(N338), .A1(N352), .B0(N672), .B1(N337), .Y(N960) );
  AOI22X1TF U610 ( .A0(N338), .A1(N349), .B0(N674), .B1(N337), .Y(N962) );
  AOI22X1TF U611 ( .A0(N335), .A1(N349), .B0(N690), .B1(N334), .Y(N970) );
  AOI22X1TF U612 ( .A0(N338), .A1(N350), .B0(N673), .B1(N337), .Y(N961) );
  AOI22X1TF U613 ( .A0(N338), .A1(N343), .B0(N671), .B1(N337), .Y(N959) );
  AOI22X1TF U614 ( .A0(N335), .A1(N346), .B0(N693), .B1(N334), .Y(N973) );
  AOI22X1TF U615 ( .A0(N340), .A1(N349), .B0(N658), .B1(N339), .Y(N954) );
  AOI22X1TF U616 ( .A0(N340), .A1(N347), .B0(N660), .B1(N339), .Y(N956) );
  AOI22X1TF U617 ( .A0(N335), .A1(N343), .B0(N687), .B1(N334), .Y(N967) );
  AOI22X1TF U618 ( .A0(N340), .A1(N346), .B0(N661), .B1(N339), .Y(N957) );
  AOI22X1TF U619 ( .A0(N335), .A1(N350), .B0(N689), .B1(N334), .Y(N969) );
  AOI22X1TF U620 ( .A0(N344), .A1(N352), .B0(N640), .B1(N342), .Y(N944) );
  AOI22X1TF U621 ( .A0(N344), .A1(N348), .B0(N643), .B1(N342), .Y(N947) );
  AOI22X1TF U622 ( .A0(N344), .A1(N350), .B0(N641), .B1(N342), .Y(N945) );
  AOI22X1TF U623 ( .A0(N353), .A1(N346), .B0(N629), .B1(N351), .Y(N941) );
  AOI22X1TF U624 ( .A0(N353), .A1(N352), .B0(N624), .B1(N351), .Y(N936) );
  AOI22X1TF U625 ( .A0(N353), .A1(N349), .B0(N626), .B1(N351), .Y(N938) );
  AOI22X1TF U626 ( .A0(N353), .A1(N350), .B0(N625), .B1(N351), .Y(N937) );
  AOI22X1TF U627 ( .A0(N353), .A1(N343), .B0(N623), .B1(N351), .Y(N1015) );
  AOI22X1TF U628 ( .A0(N353), .A1(N347), .B0(N628), .B1(N351), .Y(N940) );
  AOI22X1TF U629 ( .A0(N353), .A1(N345), .B0(N630), .B1(N351), .Y(N942) );
  AOI22X1TF U630 ( .A0(N353), .A1(N348), .B0(N627), .B1(N351), .Y(N939) );
  NAND4X2TF U631 ( .A(N22), .B(N582), .C(\OPER1_R1[2] ), .D(N336), .Y(N351) );
  AOI22X1TF U632 ( .A0(N315), .A1(N324), .B0(N684), .B1(N314), .Y(N1004) );
  AOI22X1TF U633 ( .A0(N313), .A1(N325), .B0(N699), .B1(N312), .Y(N1011) );
  AOI22X1TF U634 ( .A0(N315), .A1(N322), .B0(N686), .B1(N314), .Y(N1006) );
  AOI22X1TF U635 ( .A0(N317), .A1(N324), .B0(N668), .B1(N316), .Y(N996) );
  AOI22X1TF U636 ( .A0(N317), .A1(N330), .B0(N663), .B1(N316), .Y(N991) );
  AOI22X1TF U637 ( .A0(N313), .A1(N330), .B0(N695), .B1(N312), .Y(N1007) );
  AOI22X1TF U638 ( .A0(N315), .A1(N327), .B0(N681), .B1(N314), .Y(N1001) );
  AOI22X1TF U639 ( .A0(N315), .A1(N330), .B0(N679), .B1(N314), .Y(N999) );
  AOI22X1TF U640 ( .A0(N320), .A1(N328), .B0(N648), .B1(N319), .Y(N984) );
  AOI22X1TF U641 ( .A0(N313), .A1(N327), .B0(N697), .B1(N312), .Y(N1009) );
  AOI22X1TF U642 ( .A0(N320), .A1(N322), .B0(N654), .B1(N319), .Y(N990) );
  AOI22X1TF U643 ( .A0(N315), .A1(N325), .B0(N683), .B1(N314), .Y(N1003) );
  AOI22X1TF U644 ( .A0(N313), .A1(N324), .B0(N700), .B1(N312), .Y(N1012) );
  AOI22X1TF U645 ( .A0(N313), .A1(N322), .B0(N702), .B1(N312), .Y(N1014) );
  AOI22X1TF U646 ( .A0(N320), .A1(N327), .B0(N649), .B1(N319), .Y(N985) );
  AOI22X1TF U647 ( .A0(N317), .A1(N326), .B0(N666), .B1(N316), .Y(N994) );
  AOI22X1TF U648 ( .A0(N331), .A1(N330), .B0(N631), .B1(N329), .Y(N975) );
  AOI22X1TF U649 ( .A0(N331), .A1(N328), .B0(N632), .B1(N329), .Y(N976) );
  AOI22X1TF U650 ( .A0(N331), .A1(N322), .B0(N638), .B1(N329), .Y(N982) );
  AOI22X1TF U651 ( .A0(N331), .A1(N323), .B0(N637), .B1(N329), .Y(N981) );
  AOI22X1TF U652 ( .A0(N331), .A1(N324), .B0(N636), .B1(N329), .Y(N980) );
  AOI22X1TF U653 ( .A0(N331), .A1(N327), .B0(N633), .B1(N329), .Y(N977) );
  AOI22X1TF U654 ( .A0(N331), .A1(N325), .B0(N635), .B1(N329), .Y(N979) );
  AOI22X1TF U655 ( .A0(N331), .A1(N326), .B0(N634), .B1(N329), .Y(N978) );
  NAND4X2TF U656 ( .A(N582), .B(N22), .C(\OPER1_R1[2] ), .D(N321), .Y(N329) );
  OAI31X4TF U657 ( .A0(N1018), .A1(N308), .A2(N307), .B0(N309), .Y(N332) );
  OAI22X1TF U658 ( .A0(N935), .A1(N904), .B0(N934), .B1(N386), .Y(N307) );
  OAI211X1TF U659 ( .A0(N1204), .A1(N1185), .B0(N1145), .C0(N1144), .Y(N524)
         );
  AOI22X1TF U660 ( .A0(IO_DATAINA[12]), .A1(N206), .B0(N1215), .B1(N1160), .Y(
        N1144) );
  OAI211X1TF U661 ( .A0(N1173), .A1(N1183), .B0(N1140), .C0(N1139), .Y(N521)
         );
  AOI22X1TF U662 ( .A0(IO_DATAINB[2]), .A1(N174), .B0(D_ADDR[3]), .B1(N178), 
        .Y(N1140) );
  OAI21X1TF U663 ( .A0(N1205), .A1(N1185), .B0(N1156), .Y(N530) );
  AOI21X1TF U664 ( .A0(N206), .A1(IO_DATAINA[13]), .B0(N1155), .Y(N1156) );
  OAI22X1TF U665 ( .A0(N1204), .A1(N1183), .B0(N170), .B1(N420), .Y(N1155) );
  OAI211X1TF U666 ( .A0(N1151), .A1(N159), .B0(N1150), .C0(N1149), .Y(N527) );
  AOI22X1TF U667 ( .A0(IO_DATAINA[10]), .A1(N1202), .B0(N1213), .B1(N1206), 
        .Y(N1149) );
  OAI211X1TF U668 ( .A0(N1138), .A1(N159), .B0(N1020), .C0(N1019), .Y(N460) );
  AOI22X1TF U669 ( .A0(IO_DATAINA[3]), .A1(N1202), .B0(N1213), .B1(N1123), .Y(
        N1019) );
  AOI22X1TF U670 ( .A0(IO_DATAINB[3]), .A1(N174), .B0(D_ADDR[4]), .B1(N178), 
        .Y(N1020) );
  OAI211X1TF U671 ( .A0(N577), .A1(N814), .B0(N576), .C0(N575), .Y(N578) );
  AOI22X1TF U672 ( .A0(REG_B[2]), .A1(N574), .B0(REG_A[2]), .B1(N573), .Y(N575) );
  OAI21X1TF U673 ( .A0(REG_B[2]), .A1(N261), .B0(N728), .Y(N573) );
  AOI22X1TF U674 ( .A0(N844), .A1(N751), .B0(N502), .B1(N281), .Y(N576) );
  INVX2TF U675 ( .A(N570), .Y(N577) );
  OAI211X1TF U676 ( .A0(N246), .A1(N793), .B0(N708), .C0(N703), .Y(N570) );
  OAI22X1TF U677 ( .A0(N569), .A1(N568), .B0(N567), .B1(N853), .Y(N580) );
  OAI211X1TF U678 ( .A0(N1151), .A1(N1185), .B0(N1133), .C0(N1132), .Y(N518)
         );
  AOI22X1TF U679 ( .A0(IO_DATAINA[9]), .A1(N206), .B0(N1215), .B1(N1131), .Y(
        N1132) );
  INVX2TF U680 ( .A(N1130), .Y(N1151) );
  OAI211X1TF U681 ( .A0(N225), .A1(N621), .B0(N604), .C0(N603), .Y(N1130) );
  OAI31X1TF U682 ( .A0(N219), .A1(N829), .A2(N600), .B0(N599), .Y(N601) );
  AOI22X1TF U683 ( .A0(N846), .A1(N766), .B0(N844), .B1(N765), .Y(N599) );
  OAI211X1TF U684 ( .A0(N1209), .A1(N159), .B0(N1162), .C0(N1161), .Y(N533) );
  AOI22X1TF U685 ( .A0(IO_DATAINA[11]), .A1(N1202), .B0(N1213), .B1(N1160), 
        .Y(N1161) );
  OAI211X1TF U686 ( .A0(N227), .A1(N592), .B0(N591), .C0(N590), .Y(N1160) );
  OAI21X1TF U687 ( .A0(N849), .A1(N586), .B0(N5850), .Y(N587) );
  AOI22X1TF U688 ( .A0(N5840), .A1(N845), .B0(N846), .B1(N852), .Y(N5850) );
  INVX2TF U689 ( .A(N714), .Y(N5840) );
  OAI22X1TF U690 ( .A0(N583), .A1(N257), .B0(N727), .B1(N814), .Y(N588) );
  OAI211X1TF U691 ( .A0(N1112), .A1(N159), .B0(N1111), .C0(N1110), .Y(N5090)
         );
  AOI22X1TF U692 ( .A0(IO_DATAINA[8]), .A1(N1202), .B0(N1213), .B1(N1131), .Y(
        N1110) );
  OAI211X1TF U693 ( .A0(N224), .A1(N719), .B0(N718), .C0(N717), .Y(N1131) );
  OAI21X1TF U694 ( .A0(N714), .A1(N816), .B0(N713), .Y(N715) );
  AOI22X1TF U695 ( .A0(N846), .A1(N828), .B0(N844), .B1(N807), .Y(N713) );
  OAI22X1TF U696 ( .A0(N707), .A1(N252), .B0(N742), .B1(N814), .Y(N716) );
  INVX2TF U697 ( .A(N1109), .Y(N1112) );
  OAI211X1TF U698 ( .A0(N1173), .A1(N1185), .B0(N1172), .C0(N1171), .Y(N1174)
         );
  AOI22X1TF U699 ( .A0(N1202), .A1(IO_DATAINA[1]), .B0(N1201), .B1(
        IO_STATUS[1]), .Y(N1171) );
  AOI22X1TF U700 ( .A0(IO_DATAINB[1]), .A1(N174), .B0(D_ADDR[2]), .B1(N178), 
        .Y(N1172) );
  AOI211X1TF U701 ( .A0(REG_B[1]), .A1(N566), .B0(N565), .C0(N563), .Y(N1173)
         );
  OAI211X1TF U702 ( .A0(N561), .A1(N789), .B0(N560), .C0(N559), .Y(N563) );
  OAI211X1TF U703 ( .A0(N246), .A1(N158), .B0(N556), .C0(N555), .Y(N557) );
  OAI32X1TF U704 ( .A0(N239), .A1(REG_B[1]), .A2(N261), .B0(N728), .B1(N239), 
        .Y(N565) );
  OAI211X1TF U705 ( .A0(N1126), .A1(N159), .B0(N1105), .C0(N1104), .Y(N5060)
         );
  AOI22X1TF U706 ( .A0(IO_DATAINA[5]), .A1(N1202), .B0(N1213), .B1(N1116), .Y(
        N1104) );
  AOI22X1TF U707 ( .A0(IO_DATAINB[5]), .A1(N174), .B0(D_ADDR[6]), .B1(N1188), 
        .Y(N1105) );
  OAI211X1TF U708 ( .A0(N1126), .A1(N1185), .B0(N1125), .C0(N1124), .Y(N5150)
         );
  AOI22X1TF U709 ( .A0(IO_DATAINA[4]), .A1(N206), .B0(N1215), .B1(N1123), .Y(
        N1124) );
  AOI221X1TF U710 ( .A0(N258), .A1(N286), .B0(REG_A[3]), .B1(N203), .C0(N729), 
        .Y(N730) );
  OAI31X1TF U711 ( .A0(N789), .A1(N218), .A2(N849), .B0(N835), .Y(N729) );
  OAI21X1TF U712 ( .A0(REG_B[3]), .A1(N261), .B0(N728), .Y(N731) );
  AOI22X1TF U713 ( .A0(N844), .A1(N841), .B0(N743), .B1(N843), .Y(N733) );
  OAI211X1TF U714 ( .A0(N249), .A1(N158), .B0(N721), .C0(N720), .Y(N722) );
  AOI22X1TF U715 ( .A0(IO_DATAINB[4]), .A1(N174), .B0(D_ADDR[5]), .B1(N178), 
        .Y(N1125) );
  INVX2TF U716 ( .A(N1103), .Y(N1126) );
  OAI211X1TF U717 ( .A0(N220), .A1(N750), .B0(N749), .C0(N748), .Y(N1103) );
  OAI21X1TF U718 ( .A0(N745), .A1(N816), .B0(N744), .Y(N746) );
  AOI22X1TF U719 ( .A0(N844), .A1(N777), .B0(N743), .B1(N807), .Y(N744) );
  INVX2TF U720 ( .A(N848), .Y(N743) );
  OAI22X1TF U721 ( .A0(N741), .A1(N246), .B0(N775), .B1(N814), .Y(N747) );
  OAI211X1TF U722 ( .A0(N1119), .A1(N159), .B0(N1099), .C0(N1098), .Y(N5030)
         );
  AOI22X1TF U723 ( .A0(IO_DATAINA[7]), .A1(N206), .B0(N1213), .B1(N1109), .Y(
        N1098) );
  OAI211X1TF U724 ( .A0(N223), .A1(N856), .B0(N855), .C0(N854), .Y(N1109) );
  OAI21X1TF U725 ( .A0(N849), .A1(N848), .B0(N847), .Y(N850) );
  AOI22X1TF U726 ( .A0(N846), .A1(N845), .B0(N844), .B1(N843), .Y(N847) );
  INVX2TF U727 ( .A(N727), .Y(N843) );
  OAI22X1TF U728 ( .A0(N282), .A1(N241), .B0(N793), .B1(N248), .Y(N581) );
  AOI22X1TF U729 ( .A0(IO_DATAINB[7]), .A1(N174), .B0(D_ADDR[8]), .B1(N1188), 
        .Y(N1099) );
  OAI211X1TF U730 ( .A0(N1119), .A1(N1185), .B0(N1118), .C0(N1117), .Y(N5120)
         );
  AOI22X1TF U731 ( .A0(IO_DATAINA[6]), .A1(N206), .B0(N1215), .B1(N1116), .Y(
        N1117) );
  OAI211X1TF U732 ( .A0(N221), .A1(N774), .B0(N773), .C0(N772), .Y(N1116) );
  AOI211X1TF U733 ( .A0(N844), .A1(N771), .B0(N770), .C0(N769), .Y(N772) );
  OAI22X1TF U734 ( .A0(N799), .A1(N848), .B0(N798), .B1(N768), .Y(N769) );
  AOI22X1TF U735 ( .A0(IO_DATAINB[6]), .A1(N175), .B0(D_ADDR[7]), .B1(N178), 
        .Y(N1118) );
  INVX2TF U736 ( .A(N1097), .Y(N1119) );
  OAI211X1TF U737 ( .A0(N222), .A1(N762), .B0(N761), .C0(N760), .Y(N1097) );
  OAI31X1TF U738 ( .A0(N219), .A1(N789), .A2(N756), .B0(N755), .Y(N757) );
  AOI22X1TF U739 ( .A0(N846), .A1(N754), .B0(N844), .B1(N753), .Y(N755) );
  INVX2TF U740 ( .A(N586), .Y(N844) );
  OAI21X1TF U741 ( .A0(N170), .A1(N412), .B0(N1187), .Y(N542) );
  AOI21X1TF U742 ( .A0(N206), .A1(IO_DATAINA[15]), .B0(N1186), .Y(N1187) );
  OAI22X1TF U743 ( .A0(N230), .A1(N541), .B0(N538), .B1(N829), .Y(N544) );
  INVX2TF U744 ( .A(N567), .Y(N754) );
  AOI31X1TF U745 ( .A0(N711), .A1(N526), .A2(N706), .B0(N853), .Y(N547) );
  AOI32X1TF U746 ( .A0(N286), .A1(REG_A[14]), .A2(N230), .B0(N806), .B1(
        REG_A[14]), .Y(N548) );
  AOI32X1TF U747 ( .A0(N286), .A1(REG_A[0]), .A2(N20), .B0(N786), .B1(REG_A[0]), .Y(N787) );
  AOI211X1TF U748 ( .A0(REG_B[0]), .A1(N785), .B0(N784), .C0(N783), .Y(N788)
         );
  AOI31X1TF U749 ( .A0(N782), .A1(N781), .A2(N780), .B0(N814), .Y(N784) );
  INVX2TF U750 ( .A(N775), .Y(N776) );
  NOR4X1TF U751 ( .A(N740), .B(N739), .C(N738), .D(N737), .Y(N775) );
  NOR2X1TF U752 ( .A(N736), .B(N246), .Y(N738) );
  INVX2TF U753 ( .A(N742), .Y(N777) );
  NOR4BX1TF U754 ( .AN(N706), .B(N705), .C(N704), .D(N809), .Y(N742) );
  OAI32X4TF U755 ( .A0(N178), .A1(CODE_TYPE[4]), .A2(N240), .B0(N1018), .B1(
        N178), .Y(N1213) );
  INVX2TF U756 ( .A(N1209), .Y(N1206) );
  NOR2X1TF U757 ( .A(N793), .B(N248), .Y(N399) );
  NOR2X1TF U758 ( .A(N282), .B(N253), .Y(N550) );
  NOR2X1TF U759 ( .A(N197), .B(N241), .Y(N400) );
  AOI32X1TF U760 ( .A0(N286), .A1(REG_A[15]), .A2(N231), .B0(N786), .B1(
        REG_A[15]), .Y(N402) );
  OAI21X1TF U761 ( .A0(N853), .A1(N736), .B0(N728), .Y(N786) );
  OAI211X1TF U762 ( .A0(N243), .A1(N282), .B0(N393), .C0(N555), .Y(N845) );
  OAI211X1TF U763 ( .A0(N226), .A1(N517), .B0(N5140), .C0(N5110), .Y(N520) );
  NOR2X1TF U764 ( .A(N197), .B(N250), .Y(N705) );
  NOR2X1TF U765 ( .A(N282), .B(N255), .Y(N740) );
  OAI22X1TF U766 ( .A0(N567), .A1(N714), .B0(N569), .B1(N5050), .Y(N523) );
  AOI22X1TF U767 ( .A0(REG_B[2]), .A1(N529), .B0(N753), .B1(N218), .Y(N569) );
  OAI211X1TF U768 ( .A0(N282), .A1(N248), .B0(N5020), .C0(N808), .Y(N753) );
  AOI221X1TF U769 ( .A0(REG_B[0]), .A1(N247), .B0(N20), .B1(N241), .C0(
        REG_B[1]), .Y(N529) );
  OAI22X1TF U770 ( .A0(N197), .A1(N239), .B0(N793), .B1(N243), .Y(N5010) );
  NOR2X1TF U771 ( .A(N197), .B(N254), .Y(N739) );
  OAI21X1TF U772 ( .A0(N1205), .A1(N1204), .B0(N1203), .Y(N1211) );
  OAI22X1TF U773 ( .A0(N228), .A1(N831), .B0(N830), .B1(N829), .Y(N832) );
  NOR2X1TF U774 ( .A(N793), .B(N249), .Y(N737) );
  NOR2X1TF U775 ( .A(N736), .B(N252), .Y(N704) );
  INVX2TF U776 ( .A(N816), .Y(N820) );
  NOR2X1TF U777 ( .A(N218), .B(N219), .Y(N826) );
  NOR2X2TF U778 ( .A(REG_B[2]), .B(N219), .Y(N827) );
  OAI211X1TF U779 ( .A0(N239), .A1(N282), .B0(N709), .C0(N708), .Y(N828) );
  OAI211X1TF U780 ( .A0(N815), .A1(N814), .B0(N813), .C0(N812), .Y(N833) );
  NOR2X1TF U781 ( .A(N251), .B(N793), .Y(N809) );
  NOR2X1TF U782 ( .A(N282), .B(N250), .Y(N811) );
  INVX2TF U783 ( .A(N807), .Y(N815) );
  OAI211X1TF U784 ( .A0(N247), .A1(N282), .B0(N712), .C0(N711), .Y(N807) );
  INVX2TF U785 ( .A(N261), .Y(N287) );
  OAI211X1TF U786 ( .A0(N229), .A1(N803), .B0(N802), .C0(N801), .Y(N804) );
  AOI32X1TF U787 ( .A0(N286), .A1(REG_A[13]), .A2(N229), .B0(N806), .B1(
        REG_A[13]), .Y(N801) );
  INVX2TF U788 ( .A(N261), .Y(N286) );
  OAI22X1TF U789 ( .A0(N799), .A1(N814), .B0(N798), .B1(N797), .Y(N800) );
  AOI22X1TF U790 ( .A0(REG_B[2]), .A1(N767), .B0(N766), .B1(N218), .Y(N798) );
  OAI211X1TF U791 ( .A0(N256), .A1(N282), .B0(N598), .C0(N720), .Y(N766) );
  AOI221X1TF U792 ( .A0(N20), .A1(N239), .B0(REG_B[0]), .B1(N243), .C0(
        REG_B[1]), .Y(N767) );
  INVX2TF U793 ( .A(N840), .Y(N814) );
  INVX2TF U794 ( .A(N765), .Y(N799) );
  OAI21X1TF U795 ( .A0(N793), .A1(N247), .B0(N554), .Y(N765) );
  INVX2TF U796 ( .A(N293), .Y(N389) );
  NOR2X1TF U797 ( .A(N904), .B(N898), .Y(N293) );
  OAI32X1TF U798 ( .A0(N388), .A1(N935), .A2(N387), .B0(CODE_TYPE[4]), .B1(
        N388), .Y(N390) );
  NOR2X1TF U799 ( .A(N579), .B(N245), .Y(N387) );
  NOR2X1TF U800 ( .A(N242), .B(N386), .Y(N896) );
  OR2X2TF U801 ( .A(N901), .B(N394), .Y(N912) );
  INVX2TF U802 ( .A(N899), .Y(N394) );
  INVX2TF U803 ( .A(N935), .Y(N398) );
  INVX2TF U804 ( .A(N261), .Y(N285) );
  OR2X2TF U805 ( .A(N904), .B(N298), .Y(N261) );
  INVX2TF U806 ( .A(N406), .Y(N298) );
  INVX2TF U807 ( .A(N745), .Y(N846) );
  NOR2X2TF U808 ( .A(N218), .B(REG_B[3]), .Y(N818) );
  INVX2TF U809 ( .A(N829), .Y(N796) );
  NOR2X4TF U810 ( .A(REG_B[0]), .B(REG_B[1]), .Y(N710) );
  AOI211X1TF U811 ( .A0(REG_A[11]), .A1(N192), .B0(N792), .C0(N791), .Y(N795)
         );
  NOR2X1TF U812 ( .A(N251), .B(N282), .Y(N791) );
  NOR2X2TF U813 ( .A(N20), .B(N21), .Y(N593) );
  NOR2X1TF U814 ( .A(N197), .B(N253), .Y(N792) );
  OAI22X1TF U815 ( .A0(N291), .A1(N904), .B0(N934), .B1(N384), .Y(N838) );
  NAND2X2TF U816 ( .A(CODE_TYPE[3]), .B(N242), .Y(N904) );
  AOI21X1TF U817 ( .A0(N935), .A1(N23), .B0(N902), .Y(N291) );
  NOR2X1TF U818 ( .A(N23), .B(N1170), .Y(N1201) );
  INVX2TF U819 ( .A(N1017), .Y(N934) );
  OAI22X1TF U820 ( .A0(N179), .A1(N635), .B0(N207), .B1(N699), .Y(N919) );
  OAI22X1TF U821 ( .A0(N667), .A1(N185), .B0(N258), .B1(N183), .Y(N920) );
  OAI22X1TF U822 ( .A0(N180), .A1(N627), .B0(N1177), .B1(N691), .Y(N1157) );
  OAI22X1TF U823 ( .A0(N659), .A1(N184), .B0(N257), .B1(N182), .Y(N1158) );
  OAI22X1TF U824 ( .A0(N179), .A1(N629), .B0(N1177), .B1(N693), .Y(N1127) );
  OAI22X1TF U825 ( .A0(N661), .A1(N184), .B0(N250), .B1(N182), .Y(N1128) );
  OAI22X1TF U826 ( .A0(N179), .A1(N636), .B0(N1177), .B1(N700), .Y(N1036) );
  OAI22X1TF U827 ( .A0(N668), .A1(N184), .B0(N256), .B1(N182), .Y(N1037) );
  OAI22X1TF U828 ( .A0(N180), .A1(N631), .B0(N1177), .B1(N695), .Y(N1023) );
  OAI22X1TF U829 ( .A0(N663), .A1(N184), .B0(N255), .B1(N182), .Y(N1024) );
  OAI22X1TF U830 ( .A0(N180), .A1(N633), .B0(N1177), .B1(N697), .Y(N1100) );
  OAI22X1TF U831 ( .A0(N665), .A1(N184), .B0(N254), .B1(N182), .Y(N1101) );
  OAI22X1TF U832 ( .A0(N180), .A1(N628), .B0(N1177), .B1(N692), .Y(N1146) );
  OAI22X1TF U833 ( .A0(N660), .A1(N184), .B0(N251), .B1(N182), .Y(N1147) );
  OAI22X1TF U834 ( .A0(N180), .A1(N625), .B0(N1177), .B1(N689), .Y(N1152) );
  OAI22X1TF U835 ( .A0(N657), .A1(N184), .B0(N248), .B1(N182), .Y(N1153) );
  OAI22X1TF U836 ( .A0(N180), .A1(N630), .B0(N1177), .B1(N694), .Y(N1106) );
  OAI22X1TF U837 ( .A0(N662), .A1(N185), .B0(N252), .B1(N183), .Y(N1107) );
  OAI22X1TF U838 ( .A0(N179), .A1(N624), .B0(N207), .B1(N688), .Y(N1163) );
  OAI22X1TF U839 ( .A0(N656), .A1(N185), .B0(N241), .B1(N183), .Y(N1164) );
  OAI22X1TF U840 ( .A0(N179), .A1(N632), .B0(N207), .B1(N696), .Y(N1113) );
  OAI22X1TF U841 ( .A0(N664), .A1(N185), .B0(N249), .B1(N183), .Y(N1114) );
  OAI22X1TF U842 ( .A0(N179), .A1(N634), .B0(N207), .B1(N698), .Y(N1120) );
  OAI22X1TF U843 ( .A0(N666), .A1(N185), .B0(N246), .B1(N183), .Y(N1121) );
  OAI22X1TF U844 ( .A0(N179), .A1(N637), .B0(N207), .B1(N701), .Y(N1033) );
  OAI22X1TF U845 ( .A0(N669), .A1(N185), .B0(N239), .B1(N183), .Y(N1034) );
  OAI22X1TF U846 ( .A0(N180), .A1(N623), .B0(N207), .B1(N687), .Y(N1179) );
  OAI22X1TF U847 ( .A0(N655), .A1(N185), .B0(N247), .B1(N183), .Y(N1180) );
  OAI22X1TF U848 ( .A0(N179), .A1(N626), .B0(N207), .B1(N690), .Y(N1141) );
  OAI22X1TF U849 ( .A0(N658), .A1(N185), .B0(N253), .B1(N183), .Y(N1142) );
  OAI22X1TF U850 ( .A0(N180), .A1(N638), .B0(N1177), .B1(N702), .Y(N1030) );
  OAI22X1TF U851 ( .A0(N670), .A1(N184), .B0(N243), .B1(N182), .Y(N1031) );
  AOI211X1TF U852 ( .A0(N468), .A1(N188), .B0(N580), .C0(N578), .Y(N1138) );
  AOI211X1TF U853 ( .A0(N172), .A1(N794), .B0(N602), .C0(N601), .Y(N603) );
  AOI21X1TF U854 ( .A0(N287), .A1(N225), .B0(N166), .Y(N597) );
  AOI22X1TF U855 ( .A0(N509), .A1(N208), .B0(N475), .B1(N188), .Y(N604) );
  AOI221X1TF U856 ( .A0(N285), .A1(N250), .B0(N203), .B1(REG_A[9]), .C0(N177), 
        .Y(N621) );
  AOI211X1TF U857 ( .A0(N172), .A1(N589), .B0(N588), .C0(N587), .Y(N590) );
  AOI21X1TF U858 ( .A0(N287), .A1(N227), .B0(N166), .Y(N583) );
  AOI22X1TF U859 ( .A0(N511), .A1(N208), .B0(N477), .B1(N188), .Y(N591) );
  AOI221X1TF U860 ( .A0(N285), .A1(N257), .B0(N203), .B1(REG_A[11]), .C0(N177), 
        .Y(N592) );
  AOI211X1TF U861 ( .A0(N172), .A1(N819), .B0(N716), .C0(N715), .Y(N717) );
  AOI21X1TF U862 ( .A0(N287), .A1(N224), .B0(N166), .Y(N707) );
  AOI22X1TF U863 ( .A0(N508), .A1(N208), .B0(N474), .B1(N188), .Y(N718) );
  AOI221X1TF U864 ( .A0(N285), .A1(N252), .B0(N203), .B1(REG_A[8]), .C0(N177), 
        .Y(N719) );
  AOI22X1TF U865 ( .A0(N501), .A1(N281), .B0(N467), .B1(N187), .Y(N560) );
  AOI22X1TF U866 ( .A0(N172), .A1(N845), .B0(N840), .B1(N722), .Y(N734) );
  AOI22X1TF U867 ( .A0(N503), .A1(N281), .B0(N469), .B1(N187), .Y(N735) );
  AOI211X1TF U868 ( .A0(N172), .A1(N828), .B0(N747), .C0(N746), .Y(N748) );
  AOI21X1TF U869 ( .A0(N286), .A1(N220), .B0(N166), .Y(N741) );
  AOI22X1TF U870 ( .A0(N504), .A1(N208), .B0(N470), .B1(N188), .Y(N749) );
  AOI221X1TF U871 ( .A0(N286), .A1(N246), .B0(N203), .B1(REG_A[4]), .C0(N177), 
        .Y(N750) );
  AOI211X1TF U872 ( .A0(N172), .A1(N852), .B0(N851), .C0(N850), .Y(N854) );
  AOI211X1TF U873 ( .A0(REG_A[11]), .A1(N211), .B0(N792), .C0(N581), .Y(N727)
         );
  AOI21X1TF U874 ( .A0(N286), .A1(N223), .B0(N166), .Y(N842) );
  AOI22X1TF U875 ( .A0(N507), .A1(N281), .B0(N473), .B1(N188), .Y(N855) );
  AOI221X1TF U876 ( .A0(N285), .A1(N255), .B0(N203), .B1(REG_A[7]), .C0(N177), 
        .Y(N856) );
  AOI21X1TF U877 ( .A0(N287), .A1(N221), .B0(N166), .Y(N764) );
  AOI22X1TF U878 ( .A0(N505), .A1(N208), .B0(N471), .B1(N188), .Y(N773) );
  AOI221X1TF U879 ( .A0(N285), .A1(N254), .B0(N203), .B1(REG_A[5]), .C0(N177), 
        .Y(N774) );
  AOI211X1TF U880 ( .A0(N172), .A1(N759), .B0(N758), .C0(N757), .Y(N760) );
  AOI21X1TF U881 ( .A0(N287), .A1(N222), .B0(N166), .Y(N752) );
  AOI22X1TF U882 ( .A0(N506), .A1(N208), .B0(N472), .B1(N188), .Y(N761) );
  AOI221X1TF U883 ( .A0(N285), .A1(N249), .B0(N203), .B1(REG_A[6]), .C0(N177), 
        .Y(N762) );
  AOI221X1TF U884 ( .A0(N285), .A1(N241), .B0(N203), .B1(REG_A[14]), .C0(N177), 
        .Y(N541) );
  OAI31X1TF U885 ( .A0(N400), .A1(N550), .A2(N399), .B0(N172), .Y(N401) );
  AOI21X1TF U886 ( .A0(N710), .A1(N840), .B0(N165), .Y(N728) );
  AOI221X1TF U887 ( .A0(N285), .A1(N247), .B0(N203), .B1(REG_A[15]), .C0(N176), 
        .Y(N396) );
  AOI22X1TF U888 ( .A0(N710), .A1(REG_A[3]), .B0(N192), .B1(REG_A[1]), .Y(N393) );
  AOI22X1TF U889 ( .A0(N510), .A1(N281), .B0(N476), .B1(N187), .Y(N5110) );
  AOI22X1TF U890 ( .A0(REG_A[10]), .A1(N5080), .B0(N171), .B1(N535), .Y(N5140)
         );
  AOI221X1TF U891 ( .A0(N836), .A1(REG_A[10]), .B0(N286), .B1(N251), .C0(N176), 
        .Y(N517) );
  AOI22X1TF U892 ( .A0(REG_A[10]), .A1(N211), .B0(N192), .B1(REG_A[12]), .Y(
        N5020) );
  INVX2TF U893 ( .A(N710), .Y(N736) );
  AOI22X1TF U894 ( .A0(N710), .A1(REG_A[4]), .B0(N191), .B1(REG_A[2]), .Y(N709) );
  AOI221X1TF U895 ( .A0(N285), .A1(N253), .B0(N836), .B1(REG_A[12]), .C0(N176), 
        .Y(N831) );
  OAI31X1TF U896 ( .A0(N811), .A1(N810), .A2(N809), .B0(N171), .Y(N812) );
  AOI22X1TF U897 ( .A0(N512), .A1(N281), .B0(N478), .B1(N187), .Y(N813) );
  AOI22X1TF U898 ( .A0(N211), .A1(REG_A[12]), .B0(N192), .B1(REG_A[14]), .Y(
        N712) );
  AOI22X1TF U899 ( .A0(N710), .A1(REG_A[5]), .B0(N191), .B1(REG_A[3]), .Y(N598) );
  AOI221X1TF U900 ( .A0(N285), .A1(N248), .B0(N836), .B1(REG_A[13]), .C0(N176), 
        .Y(N803) );
  INVX2TF U901 ( .A(N1183), .Y(N1215) );
  NAND2X1TF U902 ( .A(OPER3_R3[1]), .B(N419), .Y(N1194) );
  NAND2X1TF U903 ( .A(OPER3_R3[0]), .B(N410), .Y(N1191) );
  OAI221XLTF U904 ( .A0(N579), .A1(NF), .B0(N240), .B1(N271), .C0(CODE_TYPE[2]), .Y(N295) );
  OAI2BB2XLTF U905 ( .B0(N795), .B1(N853), .A0N(N794), .A1N(N846), .Y(N805) );
  NAND2X1TF U906 ( .A(N796), .B(N818), .Y(N745) );
  CLKBUFX2TF U907 ( .A(N1194), .Y(N284) );
  CLKBUFX2TF U908 ( .A(N1191), .Y(N283) );
  INVX2TF U909 ( .A(N903), .Y(N923) );
  NAND2X1TF U910 ( .A(N562), .B(N1091), .Y(N372) );
  NOR4XLTF U911 ( .A(N24), .B(N924), .C(N923), .D(N310), .Y(N163) );
  NAND3X1TF U912 ( .A(I_ADDR[1]), .B(I_ADDR[2]), .C(I_ADDR[3]), .Y(N355) );
  NAND2X1TF U913 ( .A(N358), .B(I_ADDR[5]), .Y(N361) );
  NOR2BX1TF U914 ( .AN(N371), .B(N370), .Y(N164) );
  NAND2X1TF U915 ( .A(N905), .B(N245), .Y(N384) );
  NAND2X1TF U916 ( .A(N173), .B(N262), .Y(N898) );
  NOR4XLTF U917 ( .A(N564), .B(STATE[1]), .C(N263), .D(N294), .Y(N612) );
  NAND3X1TF U918 ( .A(N1029), .B(N383), .C(START), .Y(N301) );
  NAND2X1TF U919 ( .A(N167), .B(N302), .Y(N360) );
  AOI2BB2X1TF U920 ( .B0(I_ADDR[1]), .B1(N359), .A0N(N365), .A1N(I_ADDR[1]), 
        .Y(N303) );
  NAND2X1TF U921 ( .A(N364), .B(N270), .Y(N304) );
  NAND4X1TF U922 ( .A(N1188), .B(N311), .C(N377), .D(N306), .Y(N1016) );
  NAND2X1TF U923 ( .A(I_ADDR[1]), .B(I_ADDR[2]), .Y(N354) );
  NAND4X1TF U924 ( .A(N682), .B(N681), .C(N680), .D(N679), .Y(N374) );
  NAND2BX1TF U925 ( .AN(N898), .B(N579), .Y(N901) );
  NAND2X1TF U926 ( .A(N779), .B(REG_A[6]), .Y(N551) );
  NAND2X1TF U927 ( .A(REG_A[7]), .B(N211), .Y(N725) );
  NAND4X1TF U928 ( .A(N551), .B(N391), .C(N721), .D(N725), .Y(N852) );
  NAND2X1TF U929 ( .A(REG_A[10]), .B(N198), .Y(N549) );
  NAND2X1TF U930 ( .A(N593), .B(REG_A[8]), .Y(N552) );
  NAND2X1TF U931 ( .A(REG_A[9]), .B(N192), .Y(N724) );
  NAND4X1TF U932 ( .A(N549), .B(N552), .C(N392), .D(N724), .Y(N589) );
  NAND2X1TF U933 ( .A(N779), .B(REG_A[2]), .Y(N555) );
  AOI222XLTF U934 ( .A0(N852), .A1(N827), .B0(N589), .B1(N818), .C0(N845), 
        .C1(N826), .Y(N397) );
  OA22X1TF U935 ( .A0(N397), .A1(N829), .B0(N231), .B1(N396), .Y(N403) );
  AO21X1TF U936 ( .A0(N867), .A1(N407), .B0(N922), .Y(N1189) );
  NAND2X1TF U937 ( .A(N593), .B(REG_A[3]), .Y(N781) );
  NAND2X1TF U938 ( .A(N796), .B(N827), .Y(N714) );
  NAND2X1TF U939 ( .A(N779), .B(REG_A[11]), .Y(N808) );
  AO21X1TF U940 ( .A0(N226), .A1(N287), .B0(N166), .Y(N5080) );
  AO21X1TF U941 ( .A0(N171), .A1(N211), .B0(N165), .Y(N806) );
  NAND2X1TF U942 ( .A(N779), .B(REG_A[13]), .Y(N711) );
  NAND2X1TF U943 ( .A(N192), .B(REG_A[12]), .Y(N526) );
  NAND2X1TF U944 ( .A(N593), .B(REG_A[11]), .Y(N706) );
  NAND2X1TF U945 ( .A(N529), .B(N218), .Y(N756) );
  AOI222XLTF U946 ( .A0(N759), .A1(N827), .B0(N535), .B1(N818), .C0(N754), 
        .C1(N826), .Y(N538) );
  OAI221XLTF U947 ( .A0(REG_A[1]), .A1(N261), .B0(N239), .B1(N778), .C0(N835), 
        .Y(N566) );
  NAND2X1TF U948 ( .A(REG_A[9]), .B(N710), .Y(N596) );
  NAND2X1TF U949 ( .A(REG_A[7]), .B(N191), .Y(N595) );
  NAND4X1TF U950 ( .A(N553), .B(N595), .C(N552), .D(N551), .Y(N763) );
  AOI222XLTF U951 ( .A0(N771), .A1(N827), .B0(N763), .B1(N818), .C0(N765), 
        .C1(N826), .Y(N561) );
  NAND2X1TF U952 ( .A(N219), .B(N796), .Y(N768) );
  NAND2X1TF U953 ( .A(N218), .B(N767), .Y(N600) );
  AOI2BB2X1TF U954 ( .B0(N840), .B1(N557), .A0N(N768), .A1N(N600), .Y(N559) );
  NAND2X1TF U955 ( .A(N198), .B(REG_A[3]), .Y(N708) );
  NAND2X1TF U956 ( .A(N593), .B(REG_A[5]), .Y(N703) );
  NAND2X1TF U957 ( .A(N726), .B(N818), .Y(N586) );
  NAND2X1TF U958 ( .A(REG_A[7]), .B(N198), .Y(N622) );
  NAND4BX1TF U959 ( .AN(N811), .B(N572), .C(N571), .D(N622), .Y(N751) );
  OAI221XLTF U960 ( .A0(REG_A[2]), .A1(N261), .B0(N256), .B1(N778), .C0(N835), 
        .Y(N574) );
  NAND2X1TF U961 ( .A(N779), .B(REG_A[8]), .Y(N723) );
  NAND4X1TF U962 ( .A(N596), .B(N595), .C(N594), .D(N723), .Y(N794) );
  OAI2BB2XLTF U963 ( .B0(N597), .B1(N250), .A0N(N771), .A1N(N840), .Y(N602) );
  NAND2X1TF U964 ( .A(N198), .B(REG_A[4]), .Y(N720) );
  NAND4BBX1TF U965 ( .AN(N704), .BN(N737), .C(N703), .D(N622), .Y(N819) );
  NAND4BX1TF U966 ( .AN(N791), .B(N725), .C(N724), .D(N723), .Y(N841) );
  NAND2X1TF U967 ( .A(N726), .B(N827), .Y(N848) );
  AOI2BB2X1TF U968 ( .B0(REG_A[3]), .B1(N731), .A0N(N219), .A1N(N730), .Y(N732) );
  NAND4X1TF U969 ( .A(N735), .B(N734), .C(N733), .D(N732), .Y(N1123) );
  OAI2BB2XLTF U970 ( .B0(N752), .B1(N249), .A0N(N751), .A1N(N840), .Y(N758) );
  OAI2BB2XLTF U971 ( .B0(N764), .B1(N254), .A0N(N763), .A1N(N840), .Y(N770) );
  OAI221XLTF U972 ( .A0(REG_A[0]), .A1(N261), .B0(N243), .B1(N778), .C0(N835), 
        .Y(N785) );
  NAND2X1TF U973 ( .A(N779), .B(REG_A[1]), .Y(N782) );
  AO22X1TF U974 ( .A0(N500), .A1(N281), .B0(N466), .B1(N187), .Y(N783) );
  NAND2X1TF U975 ( .A(REG_B[3]), .B(N796), .Y(N797) );
  AO21X1TF U976 ( .A0(N287), .A1(N228), .B0(N806), .Y(N834) );
  AOI222XLTF U977 ( .A0(N828), .A1(N827), .B0(N826), .B1(N820), .C0(N819), 
        .C1(N818), .Y(N830) );
  OAI2BB2XLTF U978 ( .B0(N842), .B1(N255), .A0N(N841), .A1N(N840), .Y(N851) );
  NAND2X1TF U979 ( .A(N886), .B(N275), .Y(N868) );
  NAND2X1TF U980 ( .A(N886), .B(N273), .Y(N872) );
  NAND2X1TF U981 ( .A(N886), .B(N274), .Y(N884) );
  OAI2BB2XLTF U982 ( .B0(N905), .B1(N904), .A0N(N903), .A1N(N902), .Y(N907) );
  NAND2X1TF U983 ( .A(N913), .B(N415), .Y(N910) );
  OAI22X1TF U984 ( .A0(N416), .A1(N910), .B0(N926), .B1(N916), .Y(N1021) );
  NAND3X1TF U985 ( .A(N169), .B(N1017), .C(N935), .Y(N1170) );
  AO22X1TF U986 ( .A0(N1040), .A1(N273), .B0(N1039), .B1(I_DATAIN[6]), .Y(
        N4670) );
  AO22X1TF U987 ( .A0(N1040), .A1(N274), .B0(N1039), .B1(I_DATAIN[5]), .Y(
        N4680) );
  AO22X1TF U988 ( .A0(N1040), .A1(N275), .B0(N1039), .B1(I_DATAIN[4]), .Y(
        N4690) );
  AO22X1TF U989 ( .A0(N1040), .A1(OPER3_R3[2]), .B0(N1039), .B1(I_DATAIN[2]), 
        .Y(N4710) );
  AO22X1TF U990 ( .A0(N1040), .A1(OPER3_R3[1]), .B0(N1039), .B1(I_DATAIN[1]), 
        .Y(N4720) );
  AO22X1TF U991 ( .A0(N1040), .A1(OPER3_R3[0]), .B0(N1039), .B1(I_DATAIN[0]), 
        .Y(N4730) );
  AO22X1TF U992 ( .A0(N1042), .A1(CF_BUF), .B0(N1041), .B1(CF), .Y(N4740) );
  AO22X1TF U993 ( .A0(N1096), .A1(CODE_TYPE[3]), .B0(N1095), .B1(I_DATAIN[6]), 
        .Y(N493) );
  AO22X1TF U994 ( .A0(N1096), .A1(CODE_TYPE[2]), .B0(N1095), .B1(I_DATAIN[5]), 
        .Y(N494) );
  AO22X1TF U995 ( .A0(N1096), .A1(N24), .B0(N1095), .B1(I_DATAIN[4]), .Y(N495)
         );
  AO22X1TF U996 ( .A0(N1096), .A1(\OPER1_R1[2] ), .B0(N1095), .B1(I_DATAIN[2]), 
        .Y(N497) );
  AOI2BB2X1TF U997 ( .B0(N22), .B1(N1096), .A0N(N1096), .A1N(I_DATAIN[1]), .Y(
        N498) );
  AO22X1TF U998 ( .A0(N1096), .A1(N259), .B0(N1095), .B1(I_DATAIN[0]), .Y(N499) );
  AOI2BB2X1TF U999 ( .B0(IO_DATAINB[8]), .B1(N175), .A0N(N170), .A1N(N429), 
        .Y(N1111) );
  AOI2BB2X1TF U1000 ( .B0(IO_DATAINB[9]), .B1(N175), .A0N(N170), .A1N(N424), 
        .Y(N1133) );
  AOI2BB2X1TF U1001 ( .B0(IO_DATAINA[2]), .B1(N1202), .A0N(N1138), .A1N(N1185), 
        .Y(N1139) );
  AOI2BB2X1TF U1002 ( .B0(IO_DATAINB[12]), .B1(N175), .A0N(N170), .A1N(N423), 
        .Y(N1145) );
  AOI2BB2X1TF U1003 ( .B0(IO_DATAINB[10]), .B1(N175), .A0N(N170), .A1N(N421), 
        .Y(N1150) );
  AOI2BB2X1TF U1004 ( .B0(IO_DATAINB[11]), .B1(N175), .A0N(N170), .A1N(N418), 
        .Y(N1162) );
endmodule


module SCPU_SRAM_8BIT_ALU_SPI_TOP_VG ( CLK, RST_N, CTRL_MODE, CTRL_BGN, CPU_BGN, 
        LOAD_N, CTRL_SI, ADC_PI, CTRL_RDY, CTRL_SO, NXT, SCLK1, SCLK2, LAT, 
        SPI_SO );
  input [1:0] CTRL_MODE;
  input [15:0] ADC_PI;
  output [1:0] NXT;
  input CLK, RST_N, CTRL_BGN, CPU_BGN, LOAD_N, CTRL_SI;
  output CTRL_RDY, CTRL_SO, SCLK1, SCLK2, LAT, SPI_SO;
  wire   CEN_AFTER_MUX, WEN_AFTER_MUX, I_CLK, I_RST_N, I_CTRL_BGN, I_CPU_BGN,
         I_LOAD_N, I_CTRL_SI, I_CTRL_SO, I_SCLK1, I_SCLK2, I_SPI_SO,
         SCPU_CTRL_SPI_CEN, \SCPU_CTRL_SPI_IO_DATAOUTB[0] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[1] , \SCPU_CTRL_SPI_IO_DATAOUTB[2] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[3] , \SCPU_CTRL_SPI_IO_DATAOUTB[4] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[5] , \SCPU_CTRL_SPI_IO_DATAOUTB[6] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[7] , \SCPU_CTRL_SPI_IO_DATAOUTB[8] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[9] , \SCPU_CTRL_SPI_IO_DATAOUTB[10] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[11] , \SCPU_CTRL_SPI_IO_DATAOUTB[12] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[0] , \SCPU_CTRL_SPI_IO_DATAOUTA[1] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[2] , \SCPU_CTRL_SPI_IO_DATAOUTA[3] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[4] , \SCPU_CTRL_SPI_IO_DATAOUTA[5] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[6] , \SCPU_CTRL_SPI_IO_DATAOUTA[7] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[8] , \SCPU_CTRL_SPI_IO_DATAOUTA[9] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[10] , \SCPU_CTRL_SPI_IO_DATAOUTA[11] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[12] , \SCPU_CTRL_SPI_IO_CONTROL[0] ,
         \SCPU_CTRL_SPI_IO_CONTROL[1] , \SCPU_CTRL_SPI_IO_CONTROL[2] ,
         \SCPU_CTRL_SPI_IO_CONTROL[3] , \SCPU_CTRL_SPI_IO_CONTROL[4] ,
         \SCPU_CTRL_SPI_IO_CONTROL[5] , \SCPU_CTRL_SPI_IO_CONTROL[6] ,
         SCPU_CTRL_SPI_D_WE, SCPU_CTRL_SPI_IS_I_ADDR, SCPU_CTRL_SPI_CCT_N57,
         SCPU_CTRL_SPI_CCT_N56, SCPU_CTRL_SPI_CCT_N55, SCPU_CTRL_SPI_CCT_N53,
         SCPU_CTRL_SPI_CCT_N52, SCPU_CTRL_SPI_CCT_N51,
         SCPU_CTRL_SPI_CCT_IS_SHIFT, \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[3] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[5] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[7] , \SCPU_CTRL_SPI_CCT_REG_BITS[1] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[2] , \SCPU_CTRL_SPI_CCT_REG_BITS[3] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[4] , \SCPU_CTRL_SPI_CCT_REG_BITS[5] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[6] , \SCPU_CTRL_SPI_CCT_REG_BITS[7] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[8] , \SCPU_CTRL_SPI_CCT_REG_BITS[9] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[10] , \SCPU_CTRL_SPI_CCT_REG_BITS[11] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[12] , \SCPU_CTRL_SPI_CCT_REG_BITS[13] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[14] , \SCPU_CTRL_SPI_CCT_REG_BITS[15] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[16] , \SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ,
         SCPU_CTRL_SPI_PUT_N108, SCPU_CTRL_SPI_PUT_N107,
         SCPU_CTRL_SPI_PUT_N106, \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ,
         \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ,
         \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ,
         \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] , \SCPU_CTRL_SPI_PUT_SPI_STATE[0] ,
         \SCPU_CTRL_SPI_PUT_SPI_STATE[1] , \SCPU_CTRL_SPI_PUT_CNT_STATE[0] ,
         \SCPU_CTRL_SPI_PUT_CNT_STATE[1] , \SCPU_CTRL_SPI_PUT_CNT_STATE[2] ,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N78, N79, N80, N81, N82, N83, N84, N85, N86, N90, N92, N100,
         N103, N158, N164, N165, N189, N190, N191, N192, N193, N194, N195,
         N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206,
         N207, N208, N209, N210, N212, N213, N214, N215, N216, N218, N219,
         N220, N221, N222, N233, N234, N241, N274, N275, N276, N277, N279,
         N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292,
         N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303,
         N304, N305, N306, N307, N308, N309, N310, N311, N312, N313, N314,
         N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325,
         N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336,
         N337, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347,
         N348, N349, N350, N351, N352, N353, N354, N355, N356, N357, N358,
         N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, N369,
         N370, N371, N372, N373, N374, N375, N376, N377, N378, N379, N380,
         N381, N382, N383, N384, N385, N386, N387, N388, N389, N390, N391,
         N392, N393, N394, N395, N396, N397, N398, N399, N400, N401, N402,
         N403, N404, N405, N406, N407, N408, N409, N410, N411, N412, N413,
         N414, N415, N416, N417, N418, N419, N420, N421, N422, N423, N424,
         N425, N426, N427, N428, N429, N430, N431, N432, N433, N434;
  wire   [8:0] A_AFTER_MUX;
  wire   [7:0] D_AFTER_MUX;
  wire   [7:0] Q_FROM_SRAM;
  wire   [1:0] I_CTRL_MODE;
  wire   [15:0] I_ADC_PI;
  wire   [1:0] I_NXT;
  wire   [8:0] SCPU_CTRL_SPI_A_SPI;
  wire   [12:0] SCPU_CTRL_SPI_POUT;
  wire   [12:0] SCPU_CTRL_SPI_FOUT;
  wire   [9:0] SCPU_CTRL_SPI_IO_OFFSET;
  wire   [15:0] SCPU_CTRL_SPI_IO_DATAINA;
  wire   [0:0] SCPU_CTRL_SPI_IO_STATUS;
  wire   [7:0] SCPU_CTRL_SPI_D_DATAOUT;
  wire   [8:1] SCPU_CTRL_SPI_D_ADDR;
  wire   [8:0] SCPU_CTRL_SPI_I_ADDR;
  wire   [7:0] SCPU_CTRL_SPI_D_DATAIN;
  wire   [7:0] SCPU_CTRL_SPI_I_DATAIN;
  wire   [7:1] SCPU_CTRL_SPI_PUT_SRAM_REGS;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21;

  RA1SHD_IBM512X8 sram ( .Q(Q_FROM_SRAM), .A(A_AFTER_MUX), .D(D_AFTER_MUX), 
        .CLK(I_CLK), .CEN(CEN_AFTER_MUX), .WEN(WEN_AFTER_MUX) );
  PIC ipad_clk ( .IE(1'b1), .P(CLK), .Y(I_CLK) );
  PIC ipad_rst_n ( .IE(1'b1), .P(RST_N), .Y(I_RST_N) );
  PIC ipad_ctrl_mode0 ( .IE(1'b1), .P(CTRL_MODE[0]), .Y(I_CTRL_MODE[0]) );
  PIC ipad_ctrl_mode1 ( .IE(1'b1), .P(CTRL_MODE[1]), .Y(I_CTRL_MODE[1]) );
  PIC ipad_ctrl_bgn ( .IE(1'b1), .P(CTRL_BGN), .Y(I_CTRL_BGN) );
  PIC ipad_cpu_str ( .IE(1'b1), .P(CPU_BGN), .Y(I_CPU_BGN) );
  PIC ipad_load_n ( .IE(1'b1), .P(LOAD_N), .Y(I_LOAD_N) );
  PIC ipad_ctrl_si ( .IE(1'b1), .P(CTRL_SI), .Y(I_CTRL_SI) );
  PIC ipad_adc_pi0 ( .IE(1'b1), .P(ADC_PI[0]), .Y(I_ADC_PI[0]) );
  PIC ipad_adc_pi1 ( .IE(1'b1), .P(ADC_PI[1]), .Y(I_ADC_PI[1]) );
  PIC ipad_adc_pi2 ( .IE(1'b1), .P(ADC_PI[2]), .Y(I_ADC_PI[2]) );
  PIC ipad_adc_pi3 ( .IE(1'b1), .P(ADC_PI[3]), .Y(I_ADC_PI[3]) );
  PIC ipad_adc_pi4 ( .IE(1'b1), .P(ADC_PI[4]), .Y(I_ADC_PI[4]) );
  PIC ipad_adc_pi5 ( .IE(1'b1), .P(ADC_PI[5]), .Y(I_ADC_PI[5]) );
  PIC ipad_adc_pi6 ( .IE(1'b1), .P(ADC_PI[6]), .Y(I_ADC_PI[6]) );
  PIC ipad_adc_pi7 ( .IE(1'b1), .P(ADC_PI[7]), .Y(I_ADC_PI[7]) );
  PIC ipad_adc_pi8 ( .IE(1'b1), .P(ADC_PI[8]), .Y(I_ADC_PI[8]) );
  PIC ipad_adc_pi9 ( .IE(1'b1), .P(ADC_PI[9]), .Y(I_ADC_PI[9]) );
  PIC ipad_adc_pi10 ( .IE(1'b1), .P(ADC_PI[10]), .Y(I_ADC_PI[10]) );
  PIC ipad_adc_pi11 ( .IE(1'b1), .P(ADC_PI[11]), .Y(I_ADC_PI[11]) );
  PIC ipad_adc_pi12 ( .IE(1'b1), .P(ADC_PI[12]), .Y(I_ADC_PI[12]) );
  PIC ipad_adc_pi13 ( .IE(1'b1), .P(ADC_PI[13]), .Y(I_ADC_PI[13]) );
  PIC ipad_adc_pi14 ( .IE(1'b1), .P(ADC_PI[14]), .Y(I_ADC_PI[14]) );
  PIC ipad_adc_pi15 ( .IE(1'b1), .P(ADC_PI[15]), .Y(I_ADC_PI[15]) );
  POC8B opad_ctrl_rdy ( .A(N220), .P(CTRL_RDY) );
  POC8B opad_ctrl_so ( .A(I_CTRL_SO), .P(CTRL_SO) );
  POC8B opad_nxt0 ( .A(I_NXT[0]), .P(NXT[0]) );
  POC8B opad_nxt1 ( .A(I_NXT[1]), .P(NXT[1]) );
  POC8B opad_sclk1 ( .A(I_SCLK1), .P(SCLK1) );
  POC8B opad_sclk2 ( .A(I_SCLK2), .P(SCLK2) );
  POC8B opad_lat ( .A(N222), .P(LAT) );
  POC8B opad_spi_so ( .A(I_SPI_SO), .P(SPI_SO) );
  SHARE_SUPERALU_VG \scpu_ctrl_spi/ALU_01  ( .CLK(I_CLK), .RST_N(I_RST_N), .X_IN(
        {\SCPU_CTRL_SPI_IO_DATAOUTA[12] , \SCPU_CTRL_SPI_IO_DATAOUTA[11] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[10] , \SCPU_CTRL_SPI_IO_DATAOUTA[9] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[8] , \SCPU_CTRL_SPI_IO_DATAOUTA[7] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[6] , \SCPU_CTRL_SPI_IO_DATAOUTA[5] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[4] , \SCPU_CTRL_SPI_IO_DATAOUTA[3] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[2] , \SCPU_CTRL_SPI_IO_DATAOUTA[1] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[0] }), .Y_IN({
        \SCPU_CTRL_SPI_IO_DATAOUTB[12] , \SCPU_CTRL_SPI_IO_DATAOUTB[11] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[10] , \SCPU_CTRL_SPI_IO_DATAOUTB[9] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[8] , \SCPU_CTRL_SPI_IO_DATAOUTB[7] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[6] , \SCPU_CTRL_SPI_IO_DATAOUTB[5] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[4] , \SCPU_CTRL_SPI_IO_DATAOUTB[3] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[2] , \SCPU_CTRL_SPI_IO_DATAOUTB[1] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[0] }), .ALU_START(N396), .ALU_TYPE({
        \SCPU_CTRL_SPI_IO_CONTROL[4] , \SCPU_CTRL_SPI_IO_CONTROL[3] , 
        \SCPU_CTRL_SPI_IO_CONTROL[2] }), .MODE_TYPE({
        \SCPU_CTRL_SPI_IO_CONTROL[1] , \SCPU_CTRL_SPI_IO_CONTROL[0] }), 
        .OFFSET(SCPU_CTRL_SPI_IO_OFFSET), .FOUT(SCPU_CTRL_SPI_FOUT), .POUT(
        SCPU_CTRL_SPI_POUT), .ALU_IS_DONE(SCPU_CTRL_SPI_IO_STATUS[0]) );
  SERIAL_CPU_8BIT_VG \scpu_ctrl_spi/uut  ( .CLK(I_CLK), .ENABLE(1'b0), .RST_N(
        I_RST_N), .START(I_CPU_BGN), .I_DATAIN(SCPU_CTRL_SPI_I_DATAIN), 
        .D_DATAIN(SCPU_CTRL_SPI_D_DATAIN), .IS_I_ADDR(SCPU_CTRL_SPI_IS_I_ADDR), 
        .NXT(I_NXT), .I_ADDR(SCPU_CTRL_SPI_I_ADDR), .D_ADDR({
        SCPU_CTRL_SPI_D_ADDR, SYNOPSYS_UNCONNECTED__0}), .D_WE(
        SCPU_CTRL_SPI_D_WE), .D_DATAOUT(SCPU_CTRL_SPI_D_DATAOUT), .IO_STATUS({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, N221, SCPU_CTRL_SPI_IO_STATUS[0]}), .IO_CONTROL({
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, \SCPU_CTRL_SPI_IO_CONTROL[6] , 
        \SCPU_CTRL_SPI_IO_CONTROL[5] , \SCPU_CTRL_SPI_IO_CONTROL[4] , 
        \SCPU_CTRL_SPI_IO_CONTROL[3] , \SCPU_CTRL_SPI_IO_CONTROL[2] , 
        \SCPU_CTRL_SPI_IO_CONTROL[1] , \SCPU_CTRL_SPI_IO_CONTROL[0] }), 
        .IO_DATAINA(SCPU_CTRL_SPI_IO_DATAINA), .IO_DATAINB({1'b0, 1'b0, 1'b0, 
        SCPU_CTRL_SPI_POUT}), .IO_DATAOUTA({SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        \SCPU_CTRL_SPI_IO_DATAOUTA[12] , \SCPU_CTRL_SPI_IO_DATAOUTA[11] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[10] , \SCPU_CTRL_SPI_IO_DATAOUTA[9] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[8] , \SCPU_CTRL_SPI_IO_DATAOUTA[7] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[6] , \SCPU_CTRL_SPI_IO_DATAOUTA[5] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[4] , \SCPU_CTRL_SPI_IO_DATAOUTA[3] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[2] , \SCPU_CTRL_SPI_IO_DATAOUTA[1] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[0] }), .IO_DATAOUTB({
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, \SCPU_CTRL_SPI_IO_DATAOUTB[12] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[11] , \SCPU_CTRL_SPI_IO_DATAOUTB[10] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[9] , \SCPU_CTRL_SPI_IO_DATAOUTB[8] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[7] , \SCPU_CTRL_SPI_IO_DATAOUTB[6] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[5] , \SCPU_CTRL_SPI_IO_DATAOUTB[4] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[3] , \SCPU_CTRL_SPI_IO_DATAOUTB[2] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[1] , \SCPU_CTRL_SPI_IO_DATAOUTB[0] }), 
        .IO_OFFSET({SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SCPU_CTRL_SPI_IO_OFFSET}) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[7]  ( .D(N158), .RN(
        SCPU_CTRL_SPI_CCT_N57), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[7] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[5]  ( .D(N158), .RN(
        SCPU_CTRL_SPI_CCT_N55), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[5] ), .QN(N295) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[3]  ( .D(N158), .RN(
        SCPU_CTRL_SPI_CCT_N53), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[3] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[2]  ( .D(N158), .RN(
        SCPU_CTRL_SPI_CCT_N52), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[1]  ( .D(N158), .RN(
        SCPU_CTRL_SPI_CCT_N51), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[6]  ( .D(N158), .RN(
        SCPU_CTRL_SPI_CCT_N56), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[4]  ( .D(N45), .CK(I_CLK), 
        .SN(N44), .RN(N43), .QN(N288) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[0]  ( .D(N33), .CK(I_CLK), 
        .SN(N32), .RN(N31), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .QN(N287)
         );
  DFFSX2TF \scpu_ctrl_spi/put/cnt_state_reg[0]  ( .D(SCPU_CTRL_SPI_PUT_N106), 
        .CK(I_CLK), .SN(N274), .Q(\SCPU_CTRL_SPI_PUT_CNT_STATE[0] ), .QN(N285)
         );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[3]  ( .D(N42), .CK(I_CLK), 
        .SN(N41), .RN(N40), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] ), .QN(N284)
         );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[2]  ( .D(N39), .CK(I_CLK), 
        .SN(N38), .RN(N37), .QN(N283) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[1]  ( .D(N36), .CK(I_CLK), 
        .SN(N35), .RN(N34), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ), .QN(N282)
         );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[7]  ( .D(N189), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[7] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[6]  ( .D(N190), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[6] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[5]  ( .D(N191), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[5] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[4]  ( .D(N192), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[4] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[3]  ( .D(N193), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[3] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[2]  ( .D(N194), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[2] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[1]  ( .D(N195), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[1] ) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[7]  ( .D(N204), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[7]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[6]  ( .D(N198), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[6]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[5]  ( .D(N199), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[5]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[4]  ( .D(N200), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[4]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[3]  ( .D(N201), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[3]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[2]  ( .D(N202), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[2]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[1]  ( .D(N203), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[1]) );
  DFFTRX1TF \scpu_ctrl_spi/cct/is_shift_reg  ( .D(N164), .RN(N165), .CK(I_CLK), 
        .QN(SCPU_CTRL_SPI_CCT_IS_SHIFT) );
  DFFQX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[4]  ( .D(N215), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[0]  ( .D(N214), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[0]  ( .D(N197), .CK(I_CLK), .Q(
        I_SPI_SO) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[0]  ( .D(N196), .CK(I_CLK), .Q(
        I_CTRL_SO) );
  DFFRX1TF \scpu_ctrl_spi/put/spi_state_reg[0]  ( .D(N209), .CK(I_CLK), .RN(
        N274), .Q(\SCPU_CTRL_SPI_PUT_SPI_STATE[0] ) );
  DFFRXLTF \scpu_ctrl_spi/put/cnt_state_reg[2]  ( .D(SCPU_CTRL_SPI_PUT_N108), 
        .CK(I_CLK), .RN(N274), .Q(\SCPU_CTRL_SPI_PUT_CNT_STATE[2] ) );
  DFFNSRX4TF \scpu_ctrl_spi/put/spi_MUX_reg  ( .D(N213), .CKN(I_CLK), .SN(1'b1), .RN(1'b1), .Q(N306), .QN(N103) );
  DFFNSRXLTF \scpu_ctrl_spi/cct/D_WE_reg  ( .D(N218), .CKN(I_CLK), .SN(1'b1), 
        .RN(1'b1), .QN(N290) );
  DFFNSRX1TF \scpu_ctrl_spi/put/sram_addr_reg[7]  ( .D(N85), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[7]), .QN(N293) );
  DFFNSRXLTF \scpu_ctrl_spi/cct/CEN_reg  ( .D(N219), .CKN(I_CLK), .SN(1'b1), 
        .RN(1'b1), .Q(SCPU_CTRL_SPI_CEN) );
  DFFNSRXLTF \scpu_ctrl_spi/put/sram_addr_reg[8]  ( .D(N86), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[8]) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[15]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[16] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[15] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[14]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[15] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[14] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[13]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[14] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[13] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[12]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[13] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[12] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[11]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[12] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[11] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[10]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[11] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[10] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[9]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[10] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[9] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[8]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[9] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[8] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[16]  ( .D(I_CTRL_SI), .E(N241), 
        .CK(I_CLK), .Q(\SCPU_CTRL_SPI_CCT_REG_BITS[16] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/ctrl_state_reg[0]  ( .D(N216), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ) );
  EDFFTRXLTF \scpu_ctrl_spi/cct/ctrl_state_reg[1]  ( .RN(I_CTRL_BGN), .D(1'b1), 
        .E(N234), .CK(I_CLK), .Q(N289), .QN(N92) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_state_reg[1]  ( .D(SCPU_CTRL_SPI_PUT_N107), 
        .CK(I_CLK), .SN(1'b1), .RN(\SCPU_CTRL_SPI_IO_CONTROL[6] ), .Q(
        \SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .QN(N291) );
  DFFSRX2TF \scpu_ctrl_spi/put/spi_state_reg[2]  ( .D(N212), .CK(I_CLK), .SN(
        1'b1), .RN(\SCPU_CTRL_SPI_IO_CONTROL[6] ), .Q(N292), .QN(N100) );
  DFFSRX2TF \scpu_ctrl_spi/put/spi_state_reg[1]  ( .D(N210), .CK(I_CLK), .SN(
        1'b1), .RN(\SCPU_CTRL_SPI_IO_CONTROL[6] ), .Q(
        \SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .QN(N286) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[0]  ( .D(N205), .CK(I_CLK), 
        .SN(1'b1), .RN(\SCPU_CTRL_SPI_IO_CONTROL[6] ), .Q(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .QN(N294) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[3]  ( .D(N208), .CK(I_CLK), 
        .SN(1'b1), .RN(N274), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ), .QN(
        N297) );
  DFFRX1TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[1]  ( .D(N206), .CK(I_CLK), 
        .RN(\SCPU_CTRL_SPI_IO_CONTROL[6] ), .Q(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ) );
  DFFRX1TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[2]  ( .D(N207), .CK(I_CLK), 
        .RN(\SCPU_CTRL_SPI_IO_CONTROL[6] ), .Q(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[1]  ( .D(N79), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[1]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[3]  ( .D(N81), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[3]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[5]  ( .D(N83), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[5]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[2]  ( .D(N80), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[2]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[6]  ( .D(N84), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[6]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[4]  ( .D(N82), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[4]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[0]  ( .D(N78), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[0]), .QN(N296) );
  OR2X2TF U246 ( .A(SCPU_CTRL_SPI_IS_I_ADDR), .B(I_CTRL_BGN), .Y(N386) );
  CLKBUFX2TF U247 ( .A(N428), .Y(N300) );
  CLKBUFX2TF U248 ( .A(N428), .Y(N299) );
  INVX2TF U249 ( .A(\SCPU_CTRL_SPI_IO_CONTROL[6] ), .Y(N428) );
  NOR2BX1TF U250 ( .AN(I_ADC_PI[14]), .B(N396), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[14]) );
  AO21X1TF U251 ( .A0(N282), .A1(N430), .B0(N283), .Y(N233) );
  OAI21X1TF U252 ( .A0(N432), .A1(N433), .B0(N233), .Y(N39) );
  OA21XLTF U253 ( .A0(\SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .A1(I_CTRL_MODE[0]), 
        .B0(N329), .Y(N234) );
  CLKBUFX2TF U254 ( .A(N90), .Y(N241) );
  NOR3X1TF U273 ( .A(\SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .B(N289), .C(N328), 
        .Y(N331) );
  AOI32X1TF U274 ( .A0(SCPU_CTRL_SPI_A_SPI[0]), .A1(
        \SCPU_CTRL_SPI_IO_CONTROL[6] ), .A2(N432), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[0] ), .B1(N299), .Y(N426) );
  INVX1TF U275 ( .A(N410), .Y(N413) );
  NAND2XLTF U276 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[4] ), .B(N428), .Y(N44) );
  NAND2XLTF U277 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[3] ), .B(N428), .Y(N41) );
  NOR3BX1TF U278 ( .AN(SCPU_CTRL_SPI_CCT_IS_SHIFT), .B(N289), .C(N374), .Y(N90) );
  NAND2XLTF U279 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[2] ), .B(N428), .Y(N38) );
  NAND2XLTF U280 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[1] ), .B(N428), .Y(N35) );
  NAND2XLTF U281 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[0] ), .B(N428), .Y(N32) );
  INVX2TF U282 ( .A(\SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .Y(N374) );
  NAND2XLTF U283 ( .A(N341), .B(N397), .Y(N340) );
  CLKBUFX2TF U284 ( .A(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .Y(N396) );
  NOR2X4TF U285 ( .A(SCPU_CTRL_SPI_CEN), .B(N328), .Y(N326) );
  NAND2XLTF U286 ( .A(SCPU_CTRL_SPI_A_SPI[0]), .B(SCPU_CTRL_SPI_A_SPI[1]), .Y(
        N423) );
  NOR2X1TF U287 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .B(
        \SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .Y(N348) );
  OR2X2TF U288 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ), .B(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .Y(N301) );
  INVX2TF U289 ( .A(N428), .Y(N274) );
  INVX2TF U290 ( .A(N396), .Y(N275) );
  INVX2TF U291 ( .A(N396), .Y(N276) );
  NOR3X4TF U292 ( .A(I_CTRL_BGN), .B(N299), .C(N362), .Y(N371) );
  INVX2TF U293 ( .A(I_CTRL_BGN), .Y(N277) );
  CLKBUFX2TF U294 ( .A(N241), .Y(N298) );
  NOR3X4TF U295 ( .A(N361), .B(N360), .C(N299), .Y(N372) );
  NOR3X2TF U296 ( .A(\SCPU_CTRL_SPI_PUT_CNT_STATE[0] ), .B(
        \SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .C(\SCPU_CTRL_SPI_PUT_CNT_STATE[2] ), .Y(N397) );
  INVX2TF U297 ( .A(N432), .Y(N279) );
  NOR2BX1TF U298 ( .AN(N345), .B(N431), .Y(N429) );
  INVX2TF U299 ( .A(I_CTRL_BGN), .Y(N328) );
  AOI32X1TF U300 ( .A0(N397), .A1(N100), .A2(N341), .B0(N292), .B1(N340), .Y(
        N342) );
  NOR2X1TF U301 ( .A(N349), .B(N363), .Y(N359) );
  NAND2X1TF U302 ( .A(I_CTRL_BGN), .B(N330), .Y(N338) );
  NOR2X1TF U303 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[3] ), .B(N302), .Y(N164)
         );
  AOI222XLTF U304 ( .A0(N372), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[4]), .B0(N371), 
        .B1(Q_FROM_SRAM[4]), .C0(N370), .C1(SCPU_CTRL_SPI_PUT_SRAM_REGS[5]), 
        .Y(N367) );
  AOI222XLTF U305 ( .A0(N372), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[3]), .B0(N371), 
        .B1(Q_FROM_SRAM[3]), .C0(N370), .C1(SCPU_CTRL_SPI_PUT_SRAM_REGS[4]), 
        .Y(N366) );
  AOI222XLTF U306 ( .A0(N372), .A1(I_SPI_SO), .B0(N371), .B1(Q_FROM_SRAM[0]), 
        .C0(SCPU_CTRL_SPI_PUT_SRAM_REGS[1]), .C1(N370), .Y(N373) );
  AOI222XLTF U307 ( .A0(N372), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[1]), .B0(N371), 
        .B1(Q_FROM_SRAM[1]), .C0(N370), .C1(SCPU_CTRL_SPI_PUT_SRAM_REGS[2]), 
        .Y(N364) );
  AOI222XLTF U308 ( .A0(N372), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[2]), .B0(N371), 
        .B1(Q_FROM_SRAM[2]), .C0(N370), .C1(SCPU_CTRL_SPI_PUT_SRAM_REGS[3]), 
        .Y(N365) );
  AOI222XLTF U309 ( .A0(N372), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[5]), .B0(N371), 
        .B1(Q_FROM_SRAM[5]), .C0(N370), .C1(SCPU_CTRL_SPI_PUT_SRAM_REGS[6]), 
        .Y(N368) );
  AOI222XLTF U310 ( .A0(N372), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[6]), .B0(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[7]), .B1(N370), .C0(N371), .C1(
        Q_FROM_SRAM[6]), .Y(N369) );
  NOR2X1TF U311 ( .A(N347), .B(N100), .Y(N360) );
  NAND2X1TF U312 ( .A(N325), .B(N324), .Y(A_AFTER_MUX[8]) );
  NAND2X1TF U313 ( .A(N318), .B(N317), .Y(A_AFTER_MUX[6]) );
  NAND2X1TF U314 ( .A(N314), .B(N313), .Y(A_AFTER_MUX[4]) );
  NAND2X1TF U315 ( .A(N312), .B(N311), .Y(A_AFTER_MUX[3]) );
  NAND2X1TF U316 ( .A(N339), .B(N100), .Y(N431) );
  OR2XLTF U317 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[0] ), .B(N274), .Y(N31) );
  OR2XLTF U318 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[1] ), .B(N274), .Y(N34) );
  OR2XLTF U319 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[3] ), .B(N274), .Y(N40) );
  OR2XLTF U320 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[2] ), .B(N274), .Y(N37) );
  OR2XLTF U321 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[4] ), .B(N274), .Y(N43) );
  NOR2X1TF U322 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ), .B(N303), .Y(N304)
         );
  NAND2X1TF U323 ( .A(N295), .B(N333), .Y(N303) );
  NOR2X1TF U324 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ), .B(N334), .Y(N333)
         );
  OAI2BB2XLTF U325 ( .B0(N400), .B1(N399), .A0N(
        \SCPU_CTRL_SPI_PUT_CNT_STATE[2] ), .A1N(N398), .Y(
        SCPU_CTRL_SPI_PUT_N108) );
  NOR2X1TF U326 ( .A(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ), .B(N344), .Y(N349)
         );
  NAND2X1TF U327 ( .A(N164), .B(N165), .Y(N330) );
  OR3X1TF U328 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ), .B(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ), .C(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .Y(N302) );
  NOR2X2TF U329 ( .A(N299), .B(N363), .Y(N370) );
  NOR2X1TF U330 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .B(N286), .Y(N341) );
  NAND3X1TF U331 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .B(
        \SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .C(N100), .Y(N362) );
  NOR2BX1TF U332 ( .AN(N348), .B(N100), .Y(N222) );
  AND2X2TF U333 ( .A(N326), .B(N290), .Y(N327) );
  OAI2BB1X1TF U334 ( .A0N(\SCPU_CTRL_SPI_CCT_REG_BITS[8] ), .A1N(N326), .B0(
        N305), .Y(A_AFTER_MUX[0]) );
  NAND2X1TF U335 ( .A(\SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .B(N289), .Y(N219)
         );
  NAND2X1TF U336 ( .A(N320), .B(N319), .Y(A_AFTER_MUX[7]) );
  NAND2X1TF U337 ( .A(N316), .B(N315), .Y(A_AFTER_MUX[5]) );
  NAND2X1TF U338 ( .A(N310), .B(N309), .Y(A_AFTER_MUX[2]) );
  NAND2X1TF U339 ( .A(N308), .B(N307), .Y(A_AFTER_MUX[1]) );
  NOR2X2TF U340 ( .A(N386), .B(N306), .Y(N323) );
  NOR2X2TF U341 ( .A(N306), .B(N394), .Y(N321) );
  NAND2X2TF U342 ( .A(SCPU_CTRL_SPI_IS_I_ADDR), .B(N328), .Y(N394) );
  NOR2X2TF U343 ( .A(I_CTRL_BGN), .B(N103), .Y(N322) );
  NAND2X1TF U344 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .B(N286), .Y(N343) );
  NOR2X1TF U345 ( .A(\SCPU_CTRL_SPI_PUT_CNT_STATE[0] ), .B(N397), .Y(
        SCPU_CTRL_SPI_PUT_N106) );
  AOI21X1TF U346 ( .A0(N434), .A1(N284), .B0(N288), .Y(N45) );
  OAI31X1TF U347 ( .A0(N352), .A1(N343), .A2(N345), .B0(N342), .Y(N212) );
  OAI21X1TF U348 ( .A0(N352), .A1(N351), .B0(N350), .Y(N209) );
  OAI21X1TF U349 ( .A0(N292), .A1(N399), .B0(\SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), 
        .Y(N350) );
  AOI211X1TF U350 ( .A0(N349), .A1(N292), .B0(N348), .C0(N279), .Y(N351) );
  OAI21X1TF U351 ( .A0(N333), .A1(N295), .B0(N303), .Y(SCPU_CTRL_SPI_CCT_N55)
         );
  AOI22X1TF U352 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .A1(N279), .B0(
        N432), .B1(N287), .Y(N33) );
  OAI32X1TF U353 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ), .A1(
        \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .A2(N432), .B0(N430), .B1(N282), 
        .Y(N36) );
  OAI32X1TF U354 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] ), .A1(N433), .A2(
        N432), .B0(N434), .B1(N284), .Y(N42) );
  NOR2X1TF U355 ( .A(N431), .B(N433), .Y(N434) );
  NOR2X1TF U356 ( .A(N100), .B(N352), .Y(N346) );
  AOI21X1TF U357 ( .A0(N292), .A1(N347), .B0(N397), .Y(N352) );
  INVX2TF U358 ( .A(N338), .Y(N158) );
  NOR2X1TF U359 ( .A(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .B(N431), .Y(N430)
         );
  OAI211X1TF U360 ( .A0(N359), .A1(N294), .B0(N362), .C0(N358), .Y(N205) );
  OAI22X1TF U361 ( .A0(I_CTRL_MODE[0]), .A1(N336), .B0(N335), .B1(N338), .Y(
        N215) );
  AOI21X1TF U362 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ), .A1(N334), .B0(
        N333), .Y(N335) );
  INVX2TF U363 ( .A(N164), .Y(N334) );
  AOI22X1TF U364 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ), .A1(N354), .B0(
        N355), .B1(N297), .Y(N208) );
  AOI21X1TF U365 ( .A0(N360), .A1(N344), .B0(N400), .Y(N354) );
  OAI211X1TF U366 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .A1(N358), .B0(
        N362), .C0(N357), .Y(N206) );
  OAI21X1TF U367 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .A1(N400), .B0(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .Y(N357) );
  INVX2TF U368 ( .A(N397), .Y(N399) );
  OAI31X1TF U369 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .A1(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .A2(N400), .B0(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ), .Y(N356) );
  NOR2X1TF U370 ( .A(N361), .B(N359), .Y(N400) );
  INVX2TF U371 ( .A(N353), .Y(N344) );
  NOR3X1TF U372 ( .A(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ), .B(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .C(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .Y(N353) );
  OAI21X1TF U373 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .A1(N338), .B0(
        N337), .Y(N214) );
  INVX2TF U374 ( .A(N332), .Y(N336) );
  NOR3BX1TF U375 ( .AN(N331), .B(I_LOAD_N), .C(N330), .Y(N332) );
  NOR4X1TF U376 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[7] ), .B(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ), .C(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[5] ), .D(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ), .Y(N165) );
  OAI21X1TF U377 ( .A0(N388), .A1(N385), .B0(N377), .Y(N195) );
  AOI22X1TF U378 ( .A0(N298), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[2] ), .B0(N383), 
        .B1(\SCPU_CTRL_SPI_CCT_REG_BITS[1] ), .Y(N377) );
  OAI21X1TF U379 ( .A0(N391), .A1(N385), .B0(N380), .Y(N192) );
  AOI22X1TF U380 ( .A0(N298), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[5] ), .B0(N383), 
        .B1(\SCPU_CTRL_SPI_CCT_REG_BITS[4] ), .Y(N380) );
  OAI21X1TF U381 ( .A0(N392), .A1(N385), .B0(N381), .Y(N191) );
  AOI22X1TF U382 ( .A0(N298), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[6] ), .B0(N383), 
        .B1(\SCPU_CTRL_SPI_CCT_REG_BITS[5] ), .Y(N381) );
  OAI21X1TF U383 ( .A0(N387), .A1(N385), .B0(N376), .Y(N196) );
  AOI22X1TF U384 ( .A0(N298), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[1] ), .B0(N383), 
        .B1(I_CTRL_SO), .Y(N376) );
  OAI21X1TF U385 ( .A0(N393), .A1(N385), .B0(N382), .Y(N190) );
  AOI22X1TF U386 ( .A0(N298), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[7] ), .B0(N383), 
        .B1(\SCPU_CTRL_SPI_CCT_REG_BITS[6] ), .Y(N382) );
  OAI21X1TF U387 ( .A0(N395), .A1(N385), .B0(N384), .Y(N189) );
  AOI22X1TF U388 ( .A0(N298), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[8] ), .B0(N383), 
        .B1(\SCPU_CTRL_SPI_CCT_REG_BITS[7] ), .Y(N384) );
  OAI21X1TF U389 ( .A0(N390), .A1(N385), .B0(N379), .Y(N193) );
  AOI22X1TF U390 ( .A0(N298), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[4] ), .B0(N383), 
        .B1(\SCPU_CTRL_SPI_CCT_REG_BITS[3] ), .Y(N379) );
  OAI21X1TF U391 ( .A0(N389), .A1(N385), .B0(N378), .Y(N194) );
  AOI22X1TF U392 ( .A0(N298), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[3] ), .B0(N383), 
        .B1(\SCPU_CTRL_SPI_CCT_REG_BITS[2] ), .Y(N378) );
  NOR2X2TF U393 ( .A(N375), .B(N298), .Y(N383) );
  NAND2X2TF U394 ( .A(I_CTRL_BGN), .B(N375), .Y(N385) );
  NOR3X1TF U395 ( .A(I_CTRL_MODE[1]), .B(SCPU_CTRL_SPI_CCT_IS_SHIFT), .C(N219), 
        .Y(N375) );
  INVX2TF U396 ( .A(N367), .Y(N200) );
  INVX2TF U397 ( .A(N366), .Y(N201) );
  INVX2TF U398 ( .A(N373), .Y(N197) );
  INVX2TF U399 ( .A(N364), .Y(N203) );
  INVX2TF U400 ( .A(N365), .Y(N202) );
  INVX2TF U401 ( .A(N368), .Y(N199) );
  INVX2TF U402 ( .A(N369), .Y(N198) );
  INVX2TF U403 ( .A(N360), .Y(N363) );
  INVX2TF U404 ( .A(N341), .Y(N347) );
  INVX2TF U405 ( .A(N362), .Y(N361) );
  NOR2X1TF U406 ( .A(N92), .B(\SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .Y(N220) );
  AOI32X1TF U407 ( .A0(N103), .A1(N328), .A2(SCPU_CTRL_SPI_D_WE), .B0(
        I_CTRL_BGN), .B1(N290), .Y(WEN_AFTER_MUX) );
  NOR2X1TF U408 ( .A(N389), .B(N394), .Y(SCPU_CTRL_SPI_I_DATAIN[2]) );
  NOR2X1TF U409 ( .A(N393), .B(N394), .Y(SCPU_CTRL_SPI_I_DATAIN[6]) );
  NOR2X1TF U410 ( .A(N391), .B(N394), .Y(SCPU_CTRL_SPI_I_DATAIN[4]) );
  NOR2X1TF U411 ( .A(N387), .B(N394), .Y(SCPU_CTRL_SPI_I_DATAIN[0]) );
  NOR2X1TF U412 ( .A(N392), .B(N394), .Y(SCPU_CTRL_SPI_I_DATAIN[5]) );
  NOR2X1TF U413 ( .A(N388), .B(N394), .Y(SCPU_CTRL_SPI_I_DATAIN[1]) );
  NOR2X1TF U414 ( .A(N395), .B(N394), .Y(SCPU_CTRL_SPI_I_DATAIN[7]) );
  NOR2X1TF U415 ( .A(N390), .B(N394), .Y(SCPU_CTRL_SPI_I_DATAIN[3]) );
  NOR2X1TF U416 ( .A(N395), .B(N386), .Y(SCPU_CTRL_SPI_D_DATAIN[7]) );
  INVX2TF U417 ( .A(Q_FROM_SRAM[7]), .Y(N395) );
  NOR2X1TF U418 ( .A(N393), .B(N386), .Y(SCPU_CTRL_SPI_D_DATAIN[6]) );
  INVX2TF U419 ( .A(Q_FROM_SRAM[6]), .Y(N393) );
  NOR2X1TF U420 ( .A(N387), .B(N386), .Y(SCPU_CTRL_SPI_D_DATAIN[0]) );
  INVX2TF U421 ( .A(Q_FROM_SRAM[0]), .Y(N387) );
  NOR2X1TF U422 ( .A(N388), .B(N386), .Y(SCPU_CTRL_SPI_D_DATAIN[1]) );
  INVX2TF U423 ( .A(Q_FROM_SRAM[1]), .Y(N388) );
  NOR2X1TF U424 ( .A(N389), .B(N386), .Y(SCPU_CTRL_SPI_D_DATAIN[2]) );
  INVX2TF U425 ( .A(Q_FROM_SRAM[2]), .Y(N389) );
  NOR2X1TF U426 ( .A(N392), .B(N386), .Y(SCPU_CTRL_SPI_D_DATAIN[5]) );
  INVX2TF U427 ( .A(Q_FROM_SRAM[5]), .Y(N392) );
  NOR2X1TF U428 ( .A(N390), .B(N386), .Y(SCPU_CTRL_SPI_D_DATAIN[3]) );
  INVX2TF U429 ( .A(Q_FROM_SRAM[3]), .Y(N390) );
  NOR2X1TF U430 ( .A(N391), .B(N386), .Y(SCPU_CTRL_SPI_D_DATAIN[4]) );
  INVX2TF U431 ( .A(Q_FROM_SRAM[4]), .Y(N391) );
  OAI32X1TF U432 ( .A0(N299), .A1(N339), .A2(N103), .B0(N431), .B1(N299), .Y(
        N213) );
  OAI31X1TF U433 ( .A0(SCPU_CTRL_SPI_A_SPI[3]), .A1(N427), .A2(N420), .B0(N419), .Y(N81) );
  AOI22X1TF U434 ( .A0(SCPU_CTRL_SPI_A_SPI[3]), .A1(N418), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[3] ), .B1(N300), .Y(N419) );
  AOI21X1TF U435 ( .A0(N279), .A1(N417), .B0(N300), .Y(N418) );
  OAI31X1TF U436 ( .A0(SCPU_CTRL_SPI_A_SPI[1]), .A1(N427), .A2(N296), .B0(N425), .Y(N79) );
  AOI22X1TF U437 ( .A0(SCPU_CTRL_SPI_A_SPI[1]), .A1(N424), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[1] ), .B1(N300), .Y(N425) );
  AOI21X1TF U438 ( .A0(N279), .A1(SCPU_CTRL_SPI_A_SPI[0]), .B0(N300), .Y(N424)
         );
  OAI31X1TF U439 ( .A0(SCPU_CTRL_SPI_A_SPI[5]), .A1(N427), .A2(N413), .B0(N412), .Y(N83) );
  AOI22X1TF U440 ( .A0(SCPU_CTRL_SPI_A_SPI[5]), .A1(N411), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[5] ), .B1(N299), .Y(N412) );
  AOI21X1TF U441 ( .A0(N279), .A1(N410), .B0(N300), .Y(N411) );
  OAI31X1TF U442 ( .A0(SCPU_CTRL_SPI_A_SPI[2]), .A1(N427), .A2(N423), .B0(N422), .Y(N80) );
  AOI22X1TF U443 ( .A0(SCPU_CTRL_SPI_A_SPI[2]), .A1(N421), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[2] ), .B1(N300), .Y(N422) );
  AOI31X1TF U444 ( .A0(N279), .A1(SCPU_CTRL_SPI_A_SPI[0]), .A2(
        SCPU_CTRL_SPI_A_SPI[1]), .B0(N300), .Y(N421) );
  OAI31X1TF U445 ( .A0(SCPU_CTRL_SPI_A_SPI[4]), .A1(N427), .A2(N416), .B0(N415), .Y(N82) );
  AOI22X1TF U446 ( .A0(SCPU_CTRL_SPI_A_SPI[4]), .A1(N414), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[4] ), .B1(N300), .Y(N415) );
  AOI31X1TF U447 ( .A0(N279), .A1(N417), .A2(SCPU_CTRL_SPI_A_SPI[3]), .B0(N300), .Y(N414) );
  OAI31X1TF U448 ( .A0(SCPU_CTRL_SPI_A_SPI[6]), .A1(N427), .A2(N409), .B0(N408), .Y(N84) );
  AOI22X1TF U449 ( .A0(SCPU_CTRL_SPI_A_SPI[6]), .A1(N407), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[6] ), .B1(N299), .Y(N408) );
  AOI31X1TF U450 ( .A0(N429), .A1(N410), .A2(SCPU_CTRL_SPI_A_SPI[5]), .B0(N300), .Y(N407) );
  AOI22X1TF U451 ( .A0(N323), .A1(SCPU_CTRL_SPI_D_ADDR[8]), .B0(N326), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[16] ), .Y(N324) );
  AOI22X1TF U452 ( .A0(SCPU_CTRL_SPI_A_SPI[8]), .A1(N322), .B0(N321), .B1(
        SCPU_CTRL_SPI_I_ADDR[8]), .Y(N325) );
  AOI22X1TF U453 ( .A0(N323), .A1(SCPU_CTRL_SPI_D_ADDR[7]), .B0(N326), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[15] ), .Y(N319) );
  AOI22X1TF U454 ( .A0(SCPU_CTRL_SPI_A_SPI[7]), .A1(N322), .B0(N321), .B1(
        SCPU_CTRL_SPI_I_ADDR[7]), .Y(N320) );
  AOI22X1TF U455 ( .A0(N323), .A1(SCPU_CTRL_SPI_D_ADDR[6]), .B0(N326), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[14] ), .Y(N317) );
  AOI22X1TF U456 ( .A0(SCPU_CTRL_SPI_A_SPI[6]), .A1(N322), .B0(N321), .B1(
        SCPU_CTRL_SPI_I_ADDR[6]), .Y(N318) );
  AOI22X1TF U457 ( .A0(N323), .A1(SCPU_CTRL_SPI_D_ADDR[5]), .B0(N326), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[13] ), .Y(N315) );
  AOI22X1TF U458 ( .A0(SCPU_CTRL_SPI_A_SPI[5]), .A1(N322), .B0(N321), .B1(
        SCPU_CTRL_SPI_I_ADDR[5]), .Y(N316) );
  AOI22X1TF U459 ( .A0(N323), .A1(SCPU_CTRL_SPI_D_ADDR[4]), .B0(N326), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[12] ), .Y(N313) );
  AOI22X1TF U460 ( .A0(SCPU_CTRL_SPI_A_SPI[4]), .A1(N322), .B0(N321), .B1(
        SCPU_CTRL_SPI_I_ADDR[4]), .Y(N314) );
  AOI22X1TF U461 ( .A0(N323), .A1(SCPU_CTRL_SPI_D_ADDR[3]), .B0(N326), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[11] ), .Y(N311) );
  AOI22X1TF U462 ( .A0(SCPU_CTRL_SPI_A_SPI[3]), .A1(N322), .B0(N321), .B1(
        SCPU_CTRL_SPI_I_ADDR[3]), .Y(N312) );
  AOI22X1TF U463 ( .A0(N323), .A1(SCPU_CTRL_SPI_D_ADDR[2]), .B0(N326), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[10] ), .Y(N309) );
  AOI22X1TF U464 ( .A0(SCPU_CTRL_SPI_A_SPI[2]), .A1(N322), .B0(N321), .B1(
        SCPU_CTRL_SPI_I_ADDR[2]), .Y(N310) );
  AOI22X1TF U465 ( .A0(N323), .A1(SCPU_CTRL_SPI_D_ADDR[1]), .B0(N326), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[9] ), .Y(N307) );
  AOI22X1TF U466 ( .A0(SCPU_CTRL_SPI_A_SPI[1]), .A1(N322), .B0(N321), .B1(
        SCPU_CTRL_SPI_I_ADDR[1]), .Y(N308) );
  OAI31X1TF U467 ( .A0(SCPU_CTRL_SPI_A_SPI[8]), .A1(N293), .A2(N404), .B0(N403), .Y(N86) );
  AOI22X1TF U468 ( .A0(SCPU_CTRL_SPI_A_SPI[8]), .A1(N402), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[8] ), .B1(N299), .Y(N403) );
  OAI21X1TF U469 ( .A0(SCPU_CTRL_SPI_A_SPI[7]), .A1(N427), .B0(N406), .Y(N402)
         );
  OAI21X1TF U470 ( .A0(N406), .A1(N293), .B0(N405), .Y(N85) );
  INVX2TF U471 ( .A(N420), .Y(N417) );
  OAI21X1TF U472 ( .A0(SCPU_CTRL_SPI_A_SPI[0]), .A1(N427), .B0(N426), .Y(N78)
         );
  INVX2TF U473 ( .A(N429), .Y(N432) );
  NAND2X2TF U474 ( .A(N429), .B(\SCPU_CTRL_SPI_IO_CONTROL[6] ), .Y(N427) );
  INVX2TF U475 ( .A(N343), .Y(N339) );
  NOR2X1TF U476 ( .A(N100), .B(N343), .Y(N221) );
  NOR3X1TF U477 ( .A(N103), .B(N291), .C(N285), .Y(I_SCLK1) );
  NOR3X1TF U478 ( .A(\SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .B(N103), .C(N285), 
        .Y(I_SCLK2) );
  OAI2BB1X1TF U479 ( .A0N(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .A1N(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ), .B0(N301), .Y(
        SCPU_CTRL_SPI_CCT_N51) );
  OAI2BB1X1TF U480 ( .A0N(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ), .A1N(N301), 
        .B0(N302), .Y(SCPU_CTRL_SPI_CCT_N52) );
  OAI2BB1X1TF U481 ( .A0N(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[3] ), .A1N(N302), 
        .B0(N334), .Y(SCPU_CTRL_SPI_CCT_N53) );
  AO21X1TF U482 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ), .A1(N303), .B0(
        N304), .Y(SCPU_CTRL_SPI_CCT_N56) );
  XOR2X1TF U483 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[7] ), .B(N304), .Y(
        SCPU_CTRL_SPI_CCT_N57) );
  OAI221XLTF U484 ( .A0(N103), .A1(SCPU_CTRL_SPI_A_SPI[0]), .B0(N306), .B1(
        SCPU_CTRL_SPI_I_ADDR[0]), .C0(N328), .Y(N305) );
  NOR2BX1TF U485 ( .AN(SCPU_CTRL_SPI_CEN), .B(N328), .Y(CEN_AFTER_MUX) );
  AO22X1TF U486 ( .A0(N327), .A1(I_CTRL_SO), .B0(SCPU_CTRL_SPI_D_DATAOUT[0]), 
        .B1(N328), .Y(D_AFTER_MUX[0]) );
  AO22X1TF U487 ( .A0(N327), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[1] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[1]), .B1(N328), .Y(D_AFTER_MUX[1]) );
  AO22X1TF U488 ( .A0(N327), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[2] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[2]), .B1(N277), .Y(D_AFTER_MUX[2]) );
  AO22X1TF U489 ( .A0(N327), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[3] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[3]), .B1(N277), .Y(D_AFTER_MUX[3]) );
  AO22X1TF U490 ( .A0(N327), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[4] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[4]), .B1(N277), .Y(D_AFTER_MUX[4]) );
  AO22X1TF U491 ( .A0(N327), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[5] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[5]), .B1(N277), .Y(D_AFTER_MUX[5]) );
  AO22X1TF U492 ( .A0(N327), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[6] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[6]), .B1(N277), .Y(D_AFTER_MUX[6]) );
  AO22X1TF U493 ( .A0(N327), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[7] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[7]), .B1(N277), .Y(D_AFTER_MUX[7]) );
  NAND2BX1TF U494 ( .AN(N219), .B(I_CTRL_MODE[1]), .Y(N218) );
  OAI221XLTF U495 ( .A0(\SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .A1(I_LOAD_N), 
        .B0(N374), .B1(N330), .C0(I_CTRL_BGN), .Y(N329) );
  OAI2BB2XLTF U496 ( .B0(N374), .B1(N338), .A0N(N331), .A1N(N329), .Y(N216) );
  AO21X1TF U497 ( .A0(I_CTRL_MODE[0]), .A1(I_CTRL_MODE[1]), .B0(N336), .Y(N337) );
  NAND3X1TF U498 ( .A(N283), .B(N287), .C(N282), .Y(N433) );
  NAND3BX1TF U499 ( .AN(N433), .B(N284), .C(N288), .Y(N345) );
  OAI222X1TF U500 ( .A0(N432), .A1(N352), .B0(N347), .B1(N349), .C0(N286), 
        .C1(N346), .Y(N210) );
  NAND2X1TF U501 ( .A(N353), .B(N359), .Y(N355) );
  NAND3X1TF U502 ( .A(N362), .B(N356), .C(N355), .Y(N207) );
  NAND2X1TF U503 ( .A(N359), .B(N294), .Y(N358) );
  AO22X1TF U504 ( .A0(N372), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[7]), .B0(
        Q_FROM_SRAM[7]), .B1(N371), .Y(N204) );
  AO22X1TF U505 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[0]), .B0(N276), .B1(I_ADC_PI[0]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[0]) );
  AO22X1TF U506 ( .A0(N396), .A1(SCPU_CTRL_SPI_FOUT[10]), .B0(N275), .B1(
        I_ADC_PI[10]), .Y(SCPU_CTRL_SPI_IO_DATAINA[10]) );
  AO22X1TF U507 ( .A0(N396), .A1(SCPU_CTRL_SPI_FOUT[11]), .B0(N275), .B1(
        I_ADC_PI[11]), .Y(SCPU_CTRL_SPI_IO_DATAINA[11]) );
  AO22X1TF U508 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[12]), .B0(N276), .B1(I_ADC_PI[12]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[12]) );
  NOR2BX1TF U509 ( .AN(I_ADC_PI[13]), .B(N396), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[13]) );
  NOR2BX1TF U510 ( .AN(I_ADC_PI[15]), .B(N396), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[15]) );
  AO22X1TF U511 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[1]), .B0(N275), .B1(I_ADC_PI[1]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[1]) );
  AO22X1TF U512 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[2]), .B0(N276), .B1(I_ADC_PI[2]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[2]) );
  AO22X1TF U513 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[3]), .B0(N275), .B1(I_ADC_PI[3]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[3]) );
  AO22X1TF U514 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[4]), .B0(N276), .B1(I_ADC_PI[4]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[4]) );
  AO22X1TF U515 ( .A0(N396), .A1(SCPU_CTRL_SPI_FOUT[5]), .B0(N276), .B1(
        I_ADC_PI[5]), .Y(SCPU_CTRL_SPI_IO_DATAINA[5]) );
  AO22X1TF U516 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[6]), .B0(N276), .B1(I_ADC_PI[6]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[6]) );
  AO22X1TF U517 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[7]), .B0(N275), .B1(I_ADC_PI[7]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[7]) );
  AO22X1TF U518 ( .A0(N396), .A1(SCPU_CTRL_SPI_FOUT[8]), .B0(N276), .B1(
        I_ADC_PI[8]), .Y(SCPU_CTRL_SPI_IO_DATAINA[8]) );
  AO22X1TF U519 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[9]), .B0(N276), .B1(I_ADC_PI[9]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[9]) );
  OAI2BB2XLTF U520 ( .B0(N291), .B1(N285), .A0N(N291), .A1N(
        SCPU_CTRL_SPI_PUT_N106), .Y(SCPU_CTRL_SPI_PUT_N107) );
  NAND2X1TF U521 ( .A(N285), .B(N291), .Y(N398) );
  NAND3X1TF U522 ( .A(SCPU_CTRL_SPI_A_SPI[2]), .B(SCPU_CTRL_SPI_A_SPI[0]), .C(
        SCPU_CTRL_SPI_A_SPI[1]), .Y(N420) );
  NAND2X1TF U523 ( .A(N417), .B(SCPU_CTRL_SPI_A_SPI[3]), .Y(N416) );
  NOR2BX1TF U524 ( .AN(SCPU_CTRL_SPI_A_SPI[4]), .B(N416), .Y(N410) );
  NAND2X1TF U525 ( .A(N410), .B(SCPU_CTRL_SPI_A_SPI[5]), .Y(N409) );
  NOR2BX1TF U526 ( .AN(SCPU_CTRL_SPI_A_SPI[6]), .B(N409), .Y(N401) );
  NAND2BX1TF U527 ( .AN(N427), .B(N401), .Y(N404) );
  OAI2BB1X1TF U528 ( .A0N(N429), .A1N(N401), .B0(\SCPU_CTRL_SPI_IO_CONTROL[6] ), .Y(N406) );
  AOI2BB2X1TF U529 ( .B0(\SCPU_CTRL_SPI_IO_DATAOUTA[7] ), .B1(N299), .A0N(
        SCPU_CTRL_SPI_A_SPI[7]), .A1N(N404), .Y(N405) );
endmodule

