
module SHARE_SUPERALU_VG ( CLK, RST_N, X_IN, Y_IN, ALU_START, ALU_TYPE, MODE_TYPE, 
        OFFSET, FOUT, POUT, ALU_IS_DONE );
  input [12:0] X_IN;
  input [12:0] Y_IN;
  input [2:0] ALU_TYPE;
  input [1:0] MODE_TYPE;
  input [9:0] OFFSET;
  output [12:0] FOUT;
  output [12:0] POUT;
  input CLK, RST_N, ALU_START;
  output ALU_IS_DONE;
  wire   POST_WORK, PRE_WORK, \INDEX[2] , \RSHT_BITS[3] , SIGN_Y, C152_DATA4_0,
         C152_DATA4_1, C152_DATA4_2, C152_DATA4_3, C152_DATA4_4, C152_DATA4_5,
         C152_DATA4_6, C152_DATA4_7, C152_DATA4_8, C152_DATA4_9, C152_DATA4_10,
         C152_DATA4_11, N73, N74, N90, N91, N92, N121, N122, N123, N124, N128,
         N129, N657, N658, N659, N660, N661, N662, N663, N664, N665, N666,
         N667, N668, N669, N670, N671, N672, N673, N674, N675, N676, N677,
         N678, N679, N680, N681, N682, N683, N684, N685, N686, N687, N688,
         N689, N690, N691, N692, N693, N694, N695, N696, N697, N698, N699,
         N700, N701, N702, N703, N704, N705, N706, N707, N708, N709, N710,
         N711, N712, N713, N714, N715, N716, N717, N718, N719, N720, N721,
         N722, N723, N724, N725, N726, C2_Z_11, C2_Z_10, C2_Z_9, C2_Z_8,
         C2_Z_7, C2_Z_6, C2_Z_5, C2_Z_4, C2_Z_3, C2_Z_2, C2_Z_1,
         DP_OP_333_124_4748_N57, DP_OP_333_124_4748_N43,
         DP_OP_333_124_4748_N28, DP_OP_333_124_4748_N27,
         DP_OP_333_124_4748_N26, DP_OP_333_124_4748_N25,
         DP_OP_333_124_4748_N24, DP_OP_333_124_4748_N23,
         DP_OP_333_124_4748_N22, DP_OP_333_124_4748_N21,
         DP_OP_333_124_4748_N20, DP_OP_333_124_4748_N19,
         DP_OP_333_124_4748_N18, DP_OP_333_124_4748_N12,
         DP_OP_333_124_4748_N11, DP_OP_333_124_4748_N10, DP_OP_333_124_4748_N9,
         DP_OP_333_124_4748_N8, DP_OP_333_124_4748_N7, DP_OP_333_124_4748_N6,
         DP_OP_333_124_4748_N5, DP_OP_333_124_4748_N4, DP_OP_333_124_4748_N3,
         DP_OP_333_124_4748_N2, DP_OP_333_124_4748_N1, INTADD_0_CI,
         \INTADD_0_SUM[6] , \INTADD_0_SUM[5] , \INTADD_0_SUM[4] ,
         \INTADD_0_SUM[3] , \INTADD_0_SUM[2] , \INTADD_0_SUM[1] ,
         \INTADD_0_SUM[0] , INTADD_0_N7, INTADD_0_N6, INTADD_0_N5, INTADD_0_N4,
         INTADD_0_N3, INTADD_0_N2, INTADD_0_N1, ADD_X_132_1_N13,
         ADD_X_132_1_N12, ADD_X_132_1_N11, ADD_X_132_1_N10, ADD_X_132_1_N9,
         ADD_X_132_1_N8, ADD_X_132_1_N7, ADD_X_132_1_N6, ADD_X_132_1_N5,
         ADD_X_132_1_N4, ADD_X_132_1_N3, ADD_X_132_1_N2, N1, N2, N3, N4, N5,
         N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N77, N78, N79, N80, N81, N82,
         N83, N84, N85, N86, N87, N88, N89, N93, N94, N95, N96, N97, N98, N99,
         N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N125,
         N126, N127, N130, N131, N132, N133, N134, N135, N136, N137, N138,
         N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149,
         N150, N151, N152, N153, N154, N155, N156, N157, N158, N159, N160,
         N161, N162, N163, N164, N165, N166, N167, N168, N169, N170, N171,
         N172, N173, N174, N175, N176, N177, N178, N179, N180, N181, N182,
         N183, N184, N185, N186, N187, N188, N189, N190, N191, N192, N193,
         N194, N195, N196, N197, N198, N199, N200, N201, N202, N203, N204,
         N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215,
         N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226,
         N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237,
         N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248,
         N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259,
         N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270,
         N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281,
         N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292,
         N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303,
         N304, N305, N306, N307, N308, N309, N310, N311, N312, N313, N314,
         N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325,
         N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336,
         N337, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347,
         N348, N349, N350, N351, N352, N353, N354, N355, N356, N357, N358,
         N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, N369,
         N370, N371, N372, N373, N374, N375, N376, N377, N378, N379, N380,
         N381, N382, N383, N384, N385, N386, N387, N388, N389, N390, N391,
         N392, N393, N394, N395, N396, N397, N398, N399, N400, N401, N402,
         N403, N404, N405, N406, N407, N408, N409, N410, N411, N412, N413,
         N414, N415, N416, N417, N418, N419, N420, N421, N422, N423, N424,
         N425, N426, N427, N428, N429, N430, N431, N432, N433, N434, N435,
         N436, N437, N438, N439, N440, N441, N442, N443, N444, N445, N446,
         N447, N448, N449, N450, N451, N452, N453, N454, N455, N456, N457,
         N458, N459, N460, N461, N462, N463, N464, N465, N466, N467, N468,
         N469, N470, N471, N472, N473, N474, N475, N476, N477, N478, N479,
         N480, N481, N482, N483, N484, N485, N486, N487, N488, N489, N490,
         N491, N492, N493, N494, N495, N496, N497, N498, N499, N500, N501,
         N502, N503, N504, N505, N506, N507, N508, N509, N510, N511, N512,
         N513, N514, N515, N516, N517, N518, N519, N520, N521, N522, N523,
         N524, N525, N526, N527, N528, N529, N530, N531, N532, N533, N534,
         N535, N536, N537, N538, N539, N540, N541, N542, N543, N544, N545,
         N546, N547, N548, N549, N550, N551, N552, N553, N554, N555, N556,
         N557, N558, N559, N560, N561, N562, N563, N564, N565, N566, N567,
         N568, N569, N570, N571, N572, N573, N574, N575, N576, N577, N578,
         N579, N580, N581, N582, N583, N584, N585, N586, N587, N588, N589,
         N590, N591, N592, N593, N594, N595, N596, N597, N598, N599, N600,
         N601, N602, N603, N604, N605, N606, N607, N608, N609, N610, N611,
         N612, N613, N614, N615, N616, N617, N618, N619, N620, N621, N622,
         N623, N624, N625, N626, N627, N628, N629, N630, N631, N632, N633,
         N634, N635, N636, N637, N638, N639, N640, N641, N642, N643, N644,
         N645, N646, N647, N648, N649, N650, N651, N652, N653, N654, N655,
         N656, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736,
         N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747,
         N748, N749, N750, N751, N752, N753, N754, N755, N756, N757, N758,
         N759, N760, N761, N762, N763, N764, N765, N766, N767, N768, N769,
         N770, N771, N772, N773, N774, N775, N776, N777, N778, N779, N780,
         N781, N782, N783, N784, N785, N786, N787, N788, N789, N790, N791,
         N792, N793, N794, N795, N796, N797, N798, N799, N800, N801, N802,
         N803, N804, N805, N806, N807, N808, N809, N810, N811, N812, N813,
         N814, N815, N816, N817, N818, N819, N820, N821, N822, N823, N824,
         N825, N826, N827, N828, N829, N830, N831, N832, N833, N834, N835,
         N836, N837, N838, N839, N840, N841, N842, N843, N844, N845, N846,
         N847, N848, N849, N850, N851, N852, N853, N854, N855, N856, N857,
         N858, N859, N860, N861, N862, N863, N864, N865, N866, N867, N868,
         N869, N870, N871, N872, N873, N874, N875, N876, N877, N878, N879,
         N880, N881, N882, N883, N884, N885, N886, N887, N888, N889, N890,
         N891, N892, N893, N894, N895, N896, N897, N898, N899, N900, N901,
         N902, N903, N904, N905, N906, N907, N908, N909, N910, N911, N912,
         N913, N914, N915, N916, N917, N918, N919, N920, N921, N922, N923,
         N924, N925, N926, N927, N928, N929, N930, N931, N932, N933, N934,
         N935, N936, N937, N938, N939, N940, N941, N942, N943, N944, N945,
         N946, N947, N948, N949, N950, N951, N952, N953, N954, N955, N956,
         N957, N958, N959, N960, N961, N962, N963, N964, N965, N966, N967,
         N968, N969, N970, N971, N972, N973, N974, N975, N976, N977, N978,
         N979, N980, N981, N982, N983, N984, N985, N986, N987, N988, N989,
         N990, N991, N992, N993, N994, N995, N996, N997, N998, N999, N1000,
         N1001, N1002, N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010,
         N1011, N1012, N1013, N1014, N1015, N1016, N1017, N1018;
  wire   [12:9] XTEMP;
  wire   [12:0] DIVISION_HEAD;
  wire   [8:0] DIVISION_REMA;
  wire   [12:0] OPER_A;
  wire   [12:0] OPER_B;
  wire   [12:0] SUM_AB;
  wire   [12:0] ZTEMP;
  wire   [3:2] STEP;

  XOR2X1TF \DP_OP_333_124_4748/U27  ( .A(N77), .B(C2_Z_1), .Y(
        DP_OP_333_124_4748_N28) );
  XOR2X1TF \DP_OP_333_124_4748/U26  ( .A(N77), .B(C2_Z_2), .Y(
        DP_OP_333_124_4748_N27) );
  XOR2X1TF \DP_OP_333_124_4748/U25  ( .A(N77), .B(C2_Z_3), .Y(
        DP_OP_333_124_4748_N26) );
  XOR2X1TF \DP_OP_333_124_4748/U24  ( .A(N120), .B(C2_Z_4), .Y(
        DP_OP_333_124_4748_N25) );
  XOR2X1TF \DP_OP_333_124_4748/U23  ( .A(N77), .B(C2_Z_5), .Y(
        DP_OP_333_124_4748_N24) );
  XOR2X1TF \DP_OP_333_124_4748/U22  ( .A(N120), .B(C2_Z_6), .Y(
        DP_OP_333_124_4748_N23) );
  XOR2X1TF \DP_OP_333_124_4748/U21  ( .A(N77), .B(C2_Z_7), .Y(
        DP_OP_333_124_4748_N22) );
  XOR2X1TF \DP_OP_333_124_4748/U20  ( .A(N120), .B(C2_Z_8), .Y(
        DP_OP_333_124_4748_N21) );
  XOR2X1TF \DP_OP_333_124_4748/U19  ( .A(N77), .B(C2_Z_9), .Y(
        DP_OP_333_124_4748_N20) );
  XOR2X1TF \DP_OP_333_124_4748/U18  ( .A(N120), .B(C2_Z_10), .Y(
        DP_OP_333_124_4748_N19) );
  XOR2X1TF \DP_OP_333_124_4748/U17  ( .A(N77), .B(C2_Z_11), .Y(
        DP_OP_333_124_4748_N18) );
  ADDHXLTF \DP_OP_333_124_4748/U12  ( .A(DP_OP_333_124_4748_N28), .B(
        DP_OP_333_124_4748_N12), .CO(DP_OP_333_124_4748_N11), .S(C152_DATA4_1)
         );
  ADDHXLTF \DP_OP_333_124_4748/U11  ( .A(DP_OP_333_124_4748_N27), .B(
        DP_OP_333_124_4748_N11), .CO(DP_OP_333_124_4748_N10), .S(C152_DATA4_2)
         );
  ADDHXLTF \DP_OP_333_124_4748/U10  ( .A(DP_OP_333_124_4748_N26), .B(
        DP_OP_333_124_4748_N10), .CO(DP_OP_333_124_4748_N9), .S(C152_DATA4_3)
         );
  ADDHXLTF \DP_OP_333_124_4748/U9  ( .A(DP_OP_333_124_4748_N25), .B(
        DP_OP_333_124_4748_N9), .CO(DP_OP_333_124_4748_N8), .S(C152_DATA4_4)
         );
  ADDHXLTF \DP_OP_333_124_4748/U8  ( .A(DP_OP_333_124_4748_N24), .B(
        DP_OP_333_124_4748_N8), .CO(DP_OP_333_124_4748_N7), .S(C152_DATA4_5)
         );
  ADDHXLTF \DP_OP_333_124_4748/U7  ( .A(DP_OP_333_124_4748_N23), .B(
        DP_OP_333_124_4748_N7), .CO(DP_OP_333_124_4748_N6), .S(C152_DATA4_6)
         );
  ADDHXLTF \DP_OP_333_124_4748/U6  ( .A(DP_OP_333_124_4748_N22), .B(
        DP_OP_333_124_4748_N6), .CO(DP_OP_333_124_4748_N5), .S(C152_DATA4_7)
         );
  ADDHXLTF \DP_OP_333_124_4748/U5  ( .A(DP_OP_333_124_4748_N21), .B(
        DP_OP_333_124_4748_N5), .CO(DP_OP_333_124_4748_N4), .S(C152_DATA4_8)
         );
  ADDHXLTF \DP_OP_333_124_4748/U4  ( .A(DP_OP_333_124_4748_N20), .B(
        DP_OP_333_124_4748_N4), .CO(DP_OP_333_124_4748_N3), .S(C152_DATA4_9)
         );
  ADDHXLTF \DP_OP_333_124_4748/U3  ( .A(DP_OP_333_124_4748_N19), .B(
        DP_OP_333_124_4748_N3), .CO(DP_OP_333_124_4748_N2), .S(C152_DATA4_10)
         );
  ADDHXLTF \DP_OP_333_124_4748/U2  ( .A(DP_OP_333_124_4748_N18), .B(
        DP_OP_333_124_4748_N2), .CO(DP_OP_333_124_4748_N1), .S(C152_DATA4_11)
         );
  CMPR32X2TF \intadd_0/U8  ( .A(X_IN[1]), .B(DIVISION_HEAD[5]), .C(INTADD_0_CI), .CO(INTADD_0_N7), .S(\INTADD_0_SUM[0] ) );
  CMPR32X2TF \intadd_0/U7  ( .A(X_IN[2]), .B(DIVISION_HEAD[6]), .C(INTADD_0_N7), .CO(INTADD_0_N6), .S(\INTADD_0_SUM[1] ) );
  CMPR32X2TF \intadd_0/U6  ( .A(X_IN[3]), .B(DIVISION_HEAD[7]), .C(INTADD_0_N6), .CO(INTADD_0_N5), .S(\INTADD_0_SUM[2] ) );
  CMPR32X2TF \intadd_0/U5  ( .A(X_IN[4]), .B(DIVISION_HEAD[8]), .C(INTADD_0_N5), .CO(INTADD_0_N4), .S(\INTADD_0_SUM[3] ) );
  CMPR32X2TF \intadd_0/U4  ( .A(X_IN[5]), .B(DIVISION_HEAD[9]), .C(INTADD_0_N4), .CO(INTADD_0_N3), .S(\INTADD_0_SUM[4] ) );
  CMPR32X2TF \intadd_0/U3  ( .A(X_IN[6]), .B(DIVISION_HEAD[10]), .C(
        INTADD_0_N3), .CO(INTADD_0_N2), .S(\INTADD_0_SUM[5] ) );
  CMPR32X2TF \intadd_0/U2  ( .A(X_IN[7]), .B(DIVISION_HEAD[11]), .C(
        INTADD_0_N2), .CO(INTADD_0_N1), .S(\INTADD_0_SUM[6] ) );
  DFFRX2TF \rsht_bits_reg[3]  ( .D(N704), .CK(CLK), .RN(RST_N), .Q(
        \RSHT_BITS[3] ), .QN(N188) );
  DFFRX2TF \wtemp_reg[9]  ( .D(N673), .CK(CLK), .RN(RST_N), .Q(OPER_B[9]), 
        .QN(N187) );
  DFFRX2TF \wtemp_reg[12]  ( .D(N724), .CK(CLK), .RN(RST_N), .Q(OPER_B[12]), 
        .QN(N186) );
  DFFRX2TF \index_reg[3]  ( .D(N725), .CK(CLK), .RN(RST_N), .Q(N185), .QN(N124) );
  DFFRX2TF \wtemp_reg[11]  ( .D(N671), .CK(CLK), .RN(RST_N), .Q(OPER_B[11]), 
        .QN(N184) );
  DFFRX2TF \wtemp_reg[0]  ( .D(N682), .CK(CLK), .RN(RST_N), .Q(OPER_B[0]), 
        .QN(N183) );
  DFFRX2TF \wtemp_reg[3]  ( .D(N679), .CK(CLK), .RN(RST_N), .Q(OPER_B[3]), 
        .QN(N182) );
  DFFRX2TF \wtemp_reg[1]  ( .D(N681), .CK(CLK), .RN(RST_N), .Q(OPER_B[1]), 
        .QN(N181) );
  DFFRX2TF \index_reg[1]  ( .D(N699), .CK(CLK), .RN(RST_N), .Q(N180), .QN(N128) );
  DFFRX2TF \rsht_bits_reg[0]  ( .D(N703), .CK(CLK), .RN(RST_N), .Q(N179), .QN(
        N92) );
  DFFRX2TF \ytemp_reg[0]  ( .D(N705), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[0]), .QN(N178) );
  DFFRX2TF sign_y_reg ( .D(N694), .CK(CLK), .RN(RST_N), .Q(SIGN_Y), .QN(N177)
         );
  DFFRX2TF \wtemp_reg[4]  ( .D(N678), .CK(CLK), .RN(RST_N), .Q(OPER_B[4]), 
        .QN(N176) );
  DFFRX2TF \xtemp_reg[8]  ( .D(N711), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[12]), .QN(N175) );
  DFFSX2TF pre_work_reg ( .D(N695), .CK(CLK), .SN(RST_N), .Q(PRE_WORK), .QN(
        N174) );
  DFFRX2TF \ytemp_reg[6]  ( .D(N688), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[6]), .QN(N173) );
  DFFRX2TF \ytemp_reg[10]  ( .D(N684), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[1]), .QN(N172) );
  DFFRX2TF \ytemp_reg[2]  ( .D(N692), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[2]), .QN(N171) );
  DFFRX2TF \xtemp_reg[12]  ( .D(N723), .CK(CLK), .RN(RST_N), .Q(XTEMP[12]), 
        .QN(N170) );
  DFFRX2TF \ytemp_reg[4]  ( .D(N690), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[4]), .QN(N168) );
  DFFRX2TF \ytemp_reg[9]  ( .D(N685), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[0]), .QN(N167) );
  DFFRX2TF \ytemp_reg[7]  ( .D(N687), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[7]), .QN(N166) );
  DFFRX2TF \ytemp_reg[5]  ( .D(N689), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[5]), .QN(N165) );
  DFFRX2TF \ytemp_reg[3]  ( .D(N691), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[3]), .QN(N164) );
  DFFRX2TF \step_reg[0]  ( .D(N697), .CK(CLK), .RN(RST_N), .Q(N163), .QN(N122)
         );
  DFFRX2TF SEL_SRC_reg ( .D(N720), .CK(CLK), .RN(RST_N), .Q(POST_WORK), .QN(
        N162) );
  DFFRX2TF \ytemp_reg[11]  ( .D(N683), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[2]), .QN(N161) );
  DFFRX2TF \wtemp_reg[10]  ( .D(N672), .CK(CLK), .RN(RST_N), .Q(OPER_B[10]), 
        .QN(N160) );
  DFFRX2TF \wtemp_reg[8]  ( .D(N674), .CK(CLK), .RN(RST_N), .Q(OPER_B[8]), 
        .QN(N159) );
  DFFRX2TF \ytemp_reg[1]  ( .D(N693), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[1]), .QN(N158) );
  DFFRX2TF \rsht_bits_reg[1]  ( .D(N702), .CK(CLK), .RN(RST_N), .Q(N157), .QN(
        N91) );
  DFFRX2TF \index_reg[0]  ( .D(N726), .CK(CLK), .RN(RST_N), .Q(N156), .QN(N129) );
  DFFRX2TF \wtemp_reg[2]  ( .D(N680), .CK(CLK), .RN(RST_N), .Q(OPER_B[2]), 
        .QN(N155) );
  DFFRX2TF \xtemp_reg[11]  ( .D(N708), .CK(CLK), .RN(RST_N), .Q(XTEMP[11]), 
        .QN(N154) );
  DFFRX2TF \xtemp_reg[6]  ( .D(N713), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[10]), .QN(N153) );
  DFFRX2TF \xtemp_reg[4]  ( .D(N715), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[8]), .QN(N152) );
  DFFRX2TF \xtemp_reg[0]  ( .D(N719), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[4]), .QN(N151) );
  DFFRX2TF \xtemp_reg[2]  ( .D(N717), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[6]), .QN(N150) );
  DFFRX2TF \step_reg[3]  ( .D(N721), .CK(CLK), .RN(RST_N), .Q(STEP[3]), .QN(
        N149) );
  DFFRX2TF \step_reg[1]  ( .D(N700), .CK(CLK), .RN(RST_N), .Q(N148), .QN(N121)
         );
  DFFRX2TF \ytemp_reg[12]  ( .D(N706), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[3]), .QN(N147) );
  DFFRX2TF \xtemp_reg[10]  ( .D(N709), .CK(CLK), .RN(RST_N), .Q(XTEMP[10]), 
        .QN(N146) );
  DFFRX2TF \ytemp_reg[8]  ( .D(N686), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[8]), .QN(N145) );
  DFFRX2TF \xtemp_reg[5]  ( .D(N714), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[9]), .QN(N144) );
  DFFRX2TF \xtemp_reg[3]  ( .D(N716), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[7]), .QN(N143) );
  DFFRX2TF \xtemp_reg[1]  ( .D(N718), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[5]), .QN(N142) );
  DFFRX2TF \xtemp_reg[7]  ( .D(N712), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[11]), .QN(N141) );
  DFFRX2TF \step_reg[2]  ( .D(N696), .CK(CLK), .RN(RST_N), .Q(STEP[2]), .QN(
        N140) );
  DFFRX2TF SEL_Z_reg ( .D(N670), .CK(CLK), .RN(RST_N), .Q(N169), .QN(N123) );
  ADDHX1TF \add_x_132_1/U14  ( .A(OPER_B[0]), .B(OPER_A[0]), .CO(
        ADD_X_132_1_N13), .S(SUM_AB[0]) );
  CMPR32X2TF \add_x_132_1/U4  ( .A(OPER_A[10]), .B(OPER_B[10]), .C(
        ADD_X_132_1_N4), .CO(ADD_X_132_1_N3), .S(SUM_AB[10]) );
  CMPR32X2TF \add_x_132_1/U6  ( .A(OPER_A[8]), .B(OPER_B[8]), .C(
        ADD_X_132_1_N6), .CO(ADD_X_132_1_N5), .S(SUM_AB[8]) );
  CMPR32X2TF \add_x_132_1/U10  ( .A(OPER_A[4]), .B(OPER_B[4]), .C(
        ADD_X_132_1_N10), .CO(ADD_X_132_1_N9), .S(SUM_AB[4]) );
  CMPR32X2TF \add_x_132_1/U13  ( .A(OPER_A[1]), .B(OPER_B[1]), .C(
        ADD_X_132_1_N13), .CO(ADD_X_132_1_N12), .S(SUM_AB[1]) );
  CMPR32X2TF \add_x_132_1/U5  ( .A(OPER_A[9]), .B(OPER_B[9]), .C(
        ADD_X_132_1_N5), .CO(ADD_X_132_1_N4), .S(SUM_AB[9]) );
  CMPR32X2TF \add_x_132_1/U12  ( .A(OPER_A[2]), .B(OPER_B[2]), .C(
        ADD_X_132_1_N12), .CO(ADD_X_132_1_N11), .S(SUM_AB[2]) );
  CMPR32X2TF \add_x_132_1/U11  ( .A(OPER_A[3]), .B(OPER_B[3]), .C(
        ADD_X_132_1_N11), .CO(ADD_X_132_1_N10), .S(SUM_AB[3]) );
  CMPR32X2TF \add_x_132_1/U9  ( .A(OPER_A[5]), .B(OPER_B[5]), .C(
        ADD_X_132_1_N9), .CO(ADD_X_132_1_N8), .S(SUM_AB[5]) );
  CMPR32X2TF \add_x_132_1/U3  ( .A(OPER_A[11]), .B(OPER_B[11]), .C(
        ADD_X_132_1_N3), .CO(ADD_X_132_1_N2), .S(SUM_AB[11]) );
  DFFRX1TF \rsht_bits_reg[2]  ( .D(N701), .CK(CLK), .RN(RST_N), .QN(N90) );
  DFFRX1TF \ztemp_reg[0]  ( .D(N669), .CK(CLK), .RN(RST_N), .Q(ZTEMP[0]) );
  DFFRX1TF \wtemp_reg[6]  ( .D(N676), .CK(CLK), .RN(RST_N), .Q(OPER_B[6]) );
  DFFRX1TF \ztemp_reg[6]  ( .D(N663), .CK(CLK), .RN(RST_N), .Q(ZTEMP[6]) );
  DFFRX1TF \ztemp_reg[4]  ( .D(N665), .CK(CLK), .RN(RST_N), .Q(ZTEMP[4]) );
  DFFRX1TF \ztemp_reg[2]  ( .D(N667), .CK(CLK), .RN(RST_N), .Q(ZTEMP[2]) );
  DFFRX1TF \ztemp_reg[1]  ( .D(N668), .CK(CLK), .RN(RST_N), .Q(ZTEMP[1]) );
  DFFRX1TF \ztemp_reg[5]  ( .D(N664), .CK(CLK), .RN(RST_N), .Q(ZTEMP[5]) );
  DFFRX1TF \ztemp_reg[3]  ( .D(N666), .CK(CLK), .RN(RST_N), .Q(ZTEMP[3]) );
  DFFRX1TF \ztemp_reg[7]  ( .D(N662), .CK(CLK), .RN(RST_N), .Q(ZTEMP[7]) );
  DFFRX1TF \ztemp_reg[8]  ( .D(N661), .CK(CLK), .RN(RST_N), .Q(ZTEMP[8]) );
  DFFRX1TF \ztemp_reg[9]  ( .D(N660), .CK(CLK), .RN(RST_N), .Q(ZTEMP[9]) );
  DFFRX1TF \wtemp_reg[5]  ( .D(N677), .CK(CLK), .RN(RST_N), .Q(OPER_B[5]) );
  DFFRX1TF \wtemp_reg[7]  ( .D(N675), .CK(CLK), .RN(RST_N), .Q(OPER_B[7]) );
  DFFRX1TF \ztemp_reg[10]  ( .D(N659), .CK(CLK), .RN(RST_N), .Q(ZTEMP[10]) );
  DFFRX1TF \ztemp_reg[11]  ( .D(N658), .CK(CLK), .RN(RST_N), .Q(ZTEMP[11]) );
  DFFRX1TF \ztemp_reg[12]  ( .D(N657), .CK(CLK), .RN(RST_N), .Q(ZTEMP[12]) );
  DFFRX2TF XOR_SRC_reg ( .D(N707), .CK(CLK), .RN(RST_N), .Q(N56), .QN(N73) );
  DFFRX2TF \xtemp_reg[9]  ( .D(N710), .CK(CLK), .RN(RST_N), .Q(XTEMP[9]), .QN(
        N528) );
  DFFRX2TF sign_x_reg ( .D(N722), .CK(CLK), .RN(RST_N), .Q(N964), .QN(N74) );
  DFFRX2TF \index_reg[2]  ( .D(N698), .CK(CLK), .RN(RST_N), .Q(\INDEX[2] ) );
  NAND2X1TF U3 ( .A(ALU_START), .B(N258), .Y(N599) );
  AND2X1TF U4 ( .A(N190), .B(ZTEMP[10]), .Y(POUT[10]) );
  OAI222X1TF U5 ( .A0(N86), .A1(N170), .B0(N96), .B1(N146), .C0(N80), .C1(N147), .Y(FOUT[10]) );
  AOI21X1TF U6 ( .A0(N824), .A1(N930), .B0(N847), .Y(N1) );
  NOR3X1TF U7 ( .A(OPER_A[1]), .B(N933), .C(N824), .Y(N2) );
  OAI32X1TF U8 ( .A0(N181), .A1(OPER_B[0]), .A2(N106), .B0(N934), .B1(N181), 
        .Y(N3) );
  AOI211X1TF U9 ( .A0(OPER_B[2]), .A1(N857), .B0(N2), .C0(N3), .Y(N4) );
  OAI31X1TF U10 ( .A0(N106), .A1(N183), .A2(OPER_B[1]), .B0(N823), .Y(N5) );
  AOI211X1TF U11 ( .A0(C152_DATA4_1), .A1(N104), .B0(N885), .C0(N5), .Y(N6) );
  OAI211X1TF U12 ( .A0(N825), .A1(N1), .B0(N4), .C0(N6), .Y(N681) );
  AND2X1TF U13 ( .A(N190), .B(ZTEMP[11]), .Y(POUT[11]) );
  NOR2X1TF U14 ( .A(N97), .B(N154), .Y(FOUT[11]) );
  AOI32X1TF U15 ( .A0(N106), .A1(N836), .A2(N934), .B0(N183), .B1(N836), .Y(N7) );
  AOI211X1TF U16 ( .A0(C152_DATA4_0), .A1(N104), .B0(N885), .C0(N7), .Y(N8) );
  OAI21X1TF U17 ( .A0(N847), .A1(N930), .B0(OPER_A[0]), .Y(N9) );
  OAI211X1TF U18 ( .A0(N181), .A1(N893), .B0(N8), .C0(N9), .Y(N682) );
  NOR3X1TF U19 ( .A(Y_IN[12]), .B(Y_IN[11]), .C(Y_IN[10]), .Y(N10) );
  CLKINVX1TF U20 ( .A(N442), .Y(N11) );
  AOI22X1TF U21 ( .A0(N314), .A1(N11), .B0(N100), .B1(N736), .Y(N12) );
  OAI21X1TF U22 ( .A0(X_IN[4]), .A1(N313), .B0(N84), .Y(N13) );
  OAI22X1TF U23 ( .A0(N100), .A1(N736), .B0(X_IN[6]), .B1(N729), .Y(N14) );
  AOI31X1TF U24 ( .A0(N315), .A1(N12), .A2(N13), .B0(N14), .Y(N15) );
  AOI21X1TF U25 ( .A0(N729), .A1(X_IN[6]), .B0(N15), .Y(N16) );
  OA22X1TF U26 ( .A0(N17), .A1(N16), .B0(N488), .B1(N192), .Y(N18) );
  AO21X1TF U27 ( .A0(N468), .A1(N16), .B0(Y_IN[4]), .Y(N19) );
  AOI22X1TF U28 ( .A0(N488), .A1(N192), .B0(N18), .B1(N19), .Y(N20) );
  AOI2BB2X1TF U29 ( .B0(X_IN[9]), .B1(N20), .A0N(N502), .A1N(N83), .Y(N21) );
  CLKINVX1TF U30 ( .A(N20), .Y(N22) );
  AO21X1TF U31 ( .A0(N500), .A1(N22), .B0(Y_IN[6]), .Y(N23) );
  AOI22X1TF U32 ( .A0(Y_IN[7]), .A1(N502), .B0(N21), .B1(N23), .Y(N24) );
  AOI222XLTF U33 ( .A0(N760), .A1(X_IN[11]), .B0(N760), .B1(N24), .C0(X_IN[11]), .C1(N24), .Y(N25) );
  OAI21X1TF U34 ( .A0(Y_IN[9]), .A1(N301), .B0(N25), .Y(N26) );
  OAI211X1TF U35 ( .A0(X_IN[12]), .A1(N782), .B0(N10), .C0(N26), .Y(N768) );
  CLKINVX1TF U36 ( .A(X_IN[7]), .Y(N17) );
  AND2X1TF U37 ( .A(N190), .B(ZTEMP[12]), .Y(POUT[12]) );
  NOR2X1TF U38 ( .A(N97), .B(N170), .Y(FOUT[12]) );
  AOI22X1TF U39 ( .A0(N116), .A1(ZTEMP[0]), .B0(N1011), .B1(DIVISION_HEAD[0]), 
        .Y(N27) );
  AOI32XLTF U40 ( .A0(N1009), .A1(N27), .A2(N1018), .B0(N975), .B1(N27), .Y(
        N669) );
  OAI32X1TF U41 ( .A0(N184), .A1(N935), .A2(N106), .B0(N934), .B1(N184), .Y(
        N28) );
  CLKINVX1TF U42 ( .A(OPER_A[11]), .Y(N29) );
  OAI32X1TF U43 ( .A0(N29), .A1(N933), .A2(N932), .B0(N931), .B1(N29), .Y(N30)
         );
  AOI31X1TF U44 ( .A0(N932), .A1(N930), .A2(N29), .B0(N929), .Y(N31) );
  NOR2X1TF U45 ( .A(N105), .B(OPER_B[11]), .Y(N32) );
  AOI222XLTF U46 ( .A0(C152_DATA4_11), .A1(N103), .B0(N220), .B1(N963), .C0(
        N935), .C1(N32), .Y(N33) );
  OAI211X1TF U47 ( .A0(N186), .A1(N937), .B0(N31), .C0(N33), .Y(N34) );
  OR3X1TF U48 ( .A(N28), .B(N30), .C(N34), .Y(N671) );
  NOR2X1TF U49 ( .A(N932), .B(OPER_A[11]), .Y(N35) );
  XNOR2X1TF U50 ( .A(OPER_A[12]), .B(N35), .Y(N36) );
  AOI22X1TF U51 ( .A0(N36), .A1(N930), .B0(OPER_A[12]), .B1(N847), .Y(N37) );
  OAI21X1TF U52 ( .A0(N969), .A1(N548), .B0(N132), .Y(N38) );
  XNOR2X1TF U53 ( .A(N38), .B(N77), .Y(N39) );
  XNOR2X1TF U54 ( .A(DP_OP_333_124_4748_N1), .B(N39), .Y(N40) );
  NOR2X1TF U55 ( .A(OPER_B[11]), .B(N935), .Y(N41) );
  OAI31X1TF U56 ( .A0(N105), .A1(N41), .A2(OPER_B[12]), .B0(N823), .Y(N42) );
  AOI211X1TF U57 ( .A0(N104), .A1(N40), .B0(N929), .C0(N42), .Y(N43) );
  OAI31X1TF U58 ( .A0(OPER_B[11]), .A1(N935), .A2(N910), .B0(N867), .Y(N44) );
  AOI32X1TF U59 ( .A0(N119), .A1(OPER_B[12]), .A2(N44), .B0(N217), .B1(
        OPER_B[12]), .Y(N45) );
  NAND4BX1TF U60 ( .AN(N819), .B(N37), .C(N43), .D(N45), .Y(N724) );
  OAI21X1TF U61 ( .A0(N969), .A1(N655), .B0(N201), .Y(N46) );
  CLKMX2X2TF U62 ( .A(N77), .B(DP_OP_333_124_4748_N57), .S0(N46), .Y(
        DP_OP_333_124_4748_N12) );
  XOR2X1TF U63 ( .A(DP_OP_333_124_4748_N57), .B(N46), .Y(C152_DATA4_0) );
  NOR3X1TF U64 ( .A(N909), .B(N74), .C(N906), .Y(N47) );
  NOR2X1TF U65 ( .A(N160), .B(N937), .Y(N48) );
  AOI211X1TF U66 ( .A0(N103), .A1(C152_DATA4_9), .B0(N47), .C0(N48), .Y(N49)
         );
  NOR2X1TF U67 ( .A(N933), .B(OPER_A[9]), .Y(N50) );
  AOI22X1TF U68 ( .A0(SIGN_Y), .A1(N905), .B0(N908), .B1(N50), .Y(N51) );
  OAI21X1TF U69 ( .A0(N106), .A1(N907), .B0(N934), .Y(N52) );
  OAI21X1TF U70 ( .A0(N933), .A1(N908), .B0(N931), .Y(N53) );
  AOI22X1TF U71 ( .A0(OPER_B[9]), .A1(N52), .B0(OPER_A[9]), .B1(N53), .Y(N54)
         );
  NAND3X1TF U72 ( .A(N936), .B(N907), .C(N187), .Y(N55) );
  NAND4X1TF U73 ( .A(N49), .B(N51), .C(N54), .D(N55), .Y(N673) );
  INVX2TF U74 ( .A(N940), .Y(N110) );
  NAND2X2TF U75 ( .A(SIGN_Y), .B(N964), .Y(N970) );
  AOI22X2TF U76 ( .A0(N73), .A1(DIVISION_HEAD[3]), .B0(XTEMP[12]), .B1(N56), 
        .Y(N345) );
  OAI21XLTF U77 ( .A0(N123), .A1(N951), .B0(N950), .Y(N670) );
  NAND2X1TF U78 ( .A(N772), .B(N764), .Y(N395) );
  AND2X2TF U79 ( .A(ZTEMP[4]), .B(N133), .Y(POUT[4]) );
  NOR3BX2TF U80 ( .AN(ALU_TYPE[2]), .B(ALU_TYPE[0]), .C(ALU_TYPE[1]), .Y(N258)
         );
  OA21XLTF U81 ( .A0(SUM_AB[12]), .A1(N649), .B0(N111), .Y(N135) );
  NAND2XLTF U82 ( .A(N798), .B(SUM_AB[8]), .Y(N424) );
  NAND2X1TF U83 ( .A(N928), .B(N202), .Y(N216) );
  AOI2BB1X1TF U84 ( .A0N(N962), .A1N(N961), .B0(N960), .Y(N1010) );
  CLKINVX1TF U85 ( .A(SUM_AB[4]), .Y(N389) );
  AO21X1TF U86 ( .A0(N775), .A1(N372), .B0(N821), .Y(N509) );
  CLKINVX1TF U87 ( .A(N860), .Y(N858) );
  CLKBUFX2TF U88 ( .A(N189), .Y(DP_OP_333_124_4748_N43) );
  AND2X2TF U89 ( .A(N123), .B(N241), .Y(N256) );
  AND2XLTF U90 ( .A(\INDEX[2] ), .B(N624), .Y(N310) );
  AND2X2TF U91 ( .A(N190), .B(N73), .Y(N239) );
  AND2X2TF U92 ( .A(N109), .B(N190), .Y(N240) );
  CLKINVX1TF U93 ( .A(N620), .Y(N622) );
  CLKINVX1TF U94 ( .A(N192), .Y(N199) );
  CLKINVX1TF U95 ( .A(N832), .Y(N827) );
  CLKINVX1TF U96 ( .A(Y_IN[6]), .Y(N198) );
  CLKBUFX2TF U97 ( .A(N73), .Y(N971) );
  AOI211X1TF U98 ( .A0(X_IN[3]), .A1(N745), .B0(N440), .C0(N439), .Y(N441) );
  AOI211X1TF U99 ( .A0(Y_IN[7]), .A1(N745), .B0(N786), .C0(N785), .Y(N787) );
  AOI211X1TF U100 ( .A0(X_IN[5]), .A1(N745), .B0(N458), .C0(N457), .Y(N459) );
  OA21XLTF U101 ( .A0(SUM_AB[12]), .A1(N394), .B0(N111), .Y(N505) );
  CLKINVX2TF U102 ( .A(N864), .Y(N210) );
  AOI21X1TF U103 ( .A0(N765), .A1(N305), .B0(N386), .Y(N382) );
  INVX1TF U104 ( .A(N905), .Y(N882) );
  AND2X2TF U105 ( .A(N903), .B(N921), .Y(N936) );
  INVX2TF U106 ( .A(N114), .Y(N115) );
  OAI21XLTF U107 ( .A0(N308), .A1(N628), .B0(N621), .Y(N309) );
  OAI31X1TF U108 ( .A0(N281), .A1(X_IN[11]), .A2(N547), .B0(N280), .Y(N282) );
  AOI22X1TF U109 ( .A0(X_IN[5]), .A1(N444), .B0(N78), .B1(N98), .Y(N446) );
  AOI22X1TF U110 ( .A0(X_IN[2]), .A1(N130), .B0(X_IN[3]), .B1(N805), .Y(N784)
         );
  AOI22X1TF U111 ( .A0(X_IN[12]), .A1(N805), .B0(X_IN[11]), .B1(N130), .Y(N436) );
  AOI22X1TF U112 ( .A0(Y_IN[9]), .A1(N800), .B0(X_IN[4]), .B1(N130), .Y(N801)
         );
  OAI21X1TF U113 ( .A0(N378), .A1(N745), .B0(N380), .Y(N379) );
  AOI211X2TF U114 ( .A0(N570), .A1(N940), .B0(N594), .C0(N569), .Y(N596) );
  AOI21X1TF U115 ( .A0(N642), .A1(N119), .B0(N641), .Y(N645) );
  INVX1TF U116 ( .A(N404), .Y(N405) );
  OAI31X1TF U117 ( .A0(N564), .A1(N565), .A2(N563), .B0(N119), .Y(N581) );
  AOI32XLTF U118 ( .A0(N820), .A1(N940), .A2(N821), .B0(N637), .B1(N119), .Y(
        N643) );
  AOI22X1TF U119 ( .A0(XTEMP[11]), .A1(N125), .B0(N78), .B1(N444), .Y(N353) );
  NAND3XLTF U120 ( .A(N119), .B(N822), .C(N821), .Y(N632) );
  NAND4XLTF U121 ( .A(N611), .B(N610), .C(N609), .D(N608), .Y(N612) );
  OAI31XLTF U122 ( .A0(N111), .A1(N163), .A2(N631), .B0(N630), .Y(N636) );
  OR2X2TF U123 ( .A(N386), .B(N762), .Y(N799) );
  OAI2BB2XLTF U124 ( .B0(N760), .B1(N802), .A0N(Y_IN[6]), .A1N(N800), .Y(N777)
         );
  AOI22X1TF U125 ( .A0(X_IN[2]), .A1(N800), .B0(X_IN[3]), .B1(N444), .Y(N425)
         );
  NAND3BXLTF U126 ( .AN(N381), .B(N775), .C(N638), .Y(N365) );
  INVX1TF U127 ( .A(OPER_A[1]), .Y(N825) );
  AOI22X1TF U128 ( .A0(N192), .A1(N800), .B0(Y_IN[7]), .B1(N789), .Y(N753) );
  INVX1TF U129 ( .A(OPER_A[8]), .Y(N896) );
  AOI22X1TF U130 ( .A0(Y_IN[3]), .A1(N800), .B0(DIVISION_REMA[6]), .B1(N113), 
        .Y(N740) );
  INVX1TF U131 ( .A(OPER_A[10]), .Y(N914) );
  OAI211XLTF U132 ( .A0(N969), .A1(N364), .B0(N972), .C0(N600), .Y(N366) );
  INVX1TF U133 ( .A(OPER_A[6]), .Y(N874) );
  INVX1TF U134 ( .A(OPER_A[4]), .Y(N855) );
  AOI22X1TF U135 ( .A0(X_IN[2]), .A1(N444), .B0(X_IN[1]), .B1(N800), .Y(N418)
         );
  AOI22X1TF U136 ( .A0(Y_IN[1]), .A1(N800), .B0(DIVISION_REMA[4]), .B1(N113), 
        .Y(N730) );
  AOI22X1TF U137 ( .A0(DIVISION_HEAD[2]), .A1(N113), .B0(Y_IN[8]), .B1(N800), 
        .Y(N793) );
  AOI22X1TF U138 ( .A0(DIVISION_REMA[1]), .A1(N101), .B0(ZTEMP[1]), .B1(N169), 
        .Y(N243) );
  AOI22X1TF U139 ( .A0(DIVISION_HEAD[2]), .A1(N102), .B0(ZTEMP[11]), .B1(N134), 
        .Y(N253) );
  AOI22X1TF U140 ( .A0(DIVISION_HEAD[0]), .A1(N102), .B0(ZTEMP[9]), .B1(N134), 
        .Y(N251) );
  INVX2TF U141 ( .A(N734), .Y(N89) );
  AOI22X1TF U142 ( .A0(DIVISION_REMA[3]), .A1(N102), .B0(ZTEMP[3]), .B1(N169), 
        .Y(N245) );
  AOI22X1TF U143 ( .A0(DIVISION_REMA[0]), .A1(N101), .B0(ZTEMP[0]), .B1(N169), 
        .Y(N242) );
  AOI22X1TF U144 ( .A0(DIVISION_HEAD[1]), .A1(N102), .B0(ZTEMP[10]), .B1(N134), 
        .Y(N252) );
  INVX2TF U145 ( .A(N745), .Y(N94) );
  INVX2TF U146 ( .A(DP_OP_333_124_4748_N43), .Y(N77) );
  AOI22X1TF U147 ( .A0(DIVISION_REMA[6]), .A1(N102), .B0(ZTEMP[6]), .B1(N169), 
        .Y(N248) );
  AOI22X1TF U148 ( .A0(DIVISION_REMA[2]), .A1(N101), .B0(ZTEMP[2]), .B1(N169), 
        .Y(N244) );
  AOI22X1TF U149 ( .A0(DIVISION_REMA[8]), .A1(N102), .B0(ZTEMP[8]), .B1(N169), 
        .Y(N250) );
  AOI22X1TF U150 ( .A0(DIVISION_HEAD[3]), .A1(N102), .B0(ZTEMP[12]), .B1(N134), 
        .Y(N255) );
  AOI22X1TF U151 ( .A0(DIVISION_REMA[7]), .A1(N102), .B0(ZTEMP[7]), .B1(N169), 
        .Y(N249) );
  AOI22X1TF U152 ( .A0(DIVISION_REMA[5]), .A1(N102), .B0(ZTEMP[5]), .B1(N169), 
        .Y(N247) );
  AOI22X1TF U153 ( .A0(DIVISION_REMA[4]), .A1(N102), .B0(ZTEMP[4]), .B1(N169), 
        .Y(N246) );
  OAI21XLTF U154 ( .A0(N969), .A1(N313), .B0(N201), .Y(C2_Z_1) );
  CLKAND2X2TF U155 ( .A(N646), .B(N639), .Y(N545) );
  INVX2TF U156 ( .A(N254), .Y(N101) );
  INVX2TF U157 ( .A(N811), .Y(N112) );
  INVX1TF U158 ( .A(N341), .Y(N954) );
  AND2X2TF U159 ( .A(N341), .B(N218), .Y(N940) );
  AND2X2TF U160 ( .A(N350), .B(DP_OP_333_124_4748_N57), .Y(N745) );
  AND2X2TF U161 ( .A(N383), .B(N350), .Y(N734) );
  NAND2BXLTF U162 ( .AN(DP_OP_333_124_4748_N57), .B(N969), .Y(N202) );
  OR2X2TF U163 ( .A(N169), .B(N241), .Y(N254) );
  NAND2XLTF U164 ( .A(N218), .B(N945), .Y(N533) );
  OR3X1TF U165 ( .A(PRE_WORK), .B(N605), .C(N599), .Y(N501) );
  OR2X2TF U166 ( .A(N347), .B(N599), .Y(N811) );
  CLKAND2X2TF U167 ( .A(ZTEMP[9]), .B(N133), .Y(POUT[9]) );
  CLKAND2X2TF U168 ( .A(ZTEMP[1]), .B(N133), .Y(POUT[1]) );
  CLKAND2X2TF U169 ( .A(ZTEMP[5]), .B(N133), .Y(POUT[5]) );
  CLKAND2X2TF U170 ( .A(ZTEMP[3]), .B(N133), .Y(POUT[3]) );
  CLKAND2X2TF U171 ( .A(ZTEMP[2]), .B(N133), .Y(POUT[2]) );
  CLKAND2X2TF U172 ( .A(ZTEMP[0]), .B(N190), .Y(POUT[0]) );
  CLKAND2X2TF U173 ( .A(ZTEMP[6]), .B(N190), .Y(POUT[6]) );
  CLKAND2X2TF U174 ( .A(ZTEMP[7]), .B(N190), .Y(POUT[7]) );
  INVX2TF U175 ( .A(N195), .Y(N100) );
  CLKAND2X2TF U176 ( .A(ZTEMP[8]), .B(N190), .Y(POUT[8]) );
  INVX2TF U177 ( .A(N193), .Y(N83) );
  INVX2TF U178 ( .A(N971), .Y(N109) );
  AOI22X1TF U179 ( .A0(X_IN[11]), .A1(N547), .B0(X_IN[12]), .B1(N803), .Y(N276) );
  NAND2XLTF U180 ( .A(DIVISION_HEAD[4]), .B(N258), .Y(N221) );
  INVX2TF U181 ( .A(X_IN[3]), .Y(N194) );
  INVX2TF U182 ( .A(X_IN[5]), .Y(N195) );
  INVX1TF U183 ( .A(X_IN[2]), .Y(N770) );
  INVX2TF U184 ( .A(Y_IN[7]), .Y(N193) );
  INVX2TF U185 ( .A(N297), .Y(N78) );
  INVX2TF U186 ( .A(N240), .Y(N79) );
  INVX2TF U187 ( .A(N240), .Y(N80) );
  INVX2TF U188 ( .A(N1018), .Y(N81) );
  INVX2TF U189 ( .A(N1018), .Y(N82) );
  INVX2TF U190 ( .A(N194), .Y(N84) );
  INVX2TF U191 ( .A(N239), .Y(N85) );
  INVX2TF U192 ( .A(N239), .Y(N86) );
  INVX2TF U193 ( .A(N501), .Y(N87) );
  INVX2TF U194 ( .A(N501), .Y(N88) );
  INVX2TF U195 ( .A(N734), .Y(N93) );
  INVX2TF U196 ( .A(N745), .Y(N95) );
  INVX2TF U197 ( .A(N258), .Y(N96) );
  INVX2TF U198 ( .A(N258), .Y(N97) );
  INVX2TF U199 ( .A(N395), .Y(N98) );
  INVX2TF U200 ( .A(N395), .Y(N99) );
  INVX2TF U201 ( .A(N254), .Y(N102) );
  INVX2TF U202 ( .A(N216), .Y(N103) );
  INVX2TF U203 ( .A(N216), .Y(N104) );
  INVX2TF U204 ( .A(N936), .Y(N105) );
  INVX2TF U205 ( .A(N936), .Y(N106) );
  INVX2TF U206 ( .A(N256), .Y(N107) );
  INVX2TF U207 ( .A(N256), .Y(N108) );
  INVX2TF U208 ( .A(N940), .Y(N111) );
  INVX2TF U209 ( .A(N811), .Y(N113) );
  INVX2TF U210 ( .A(N1010), .Y(N114) );
  INVX2TF U211 ( .A(N114), .Y(N116) );
  INVX2TF U212 ( .A(N509), .Y(N117) );
  INVX2TF U213 ( .A(N509), .Y(N118) );
  INVX2TF U214 ( .A(N110), .Y(N119) );
  INVX2TF U215 ( .A(DP_OP_333_124_4748_N43), .Y(N120) );
  INVX2TF U216 ( .A(N89), .Y(N125) );
  AOI222X4TF U217 ( .A0(N487), .A1(N146), .B0(N487), .B1(N502), .C0(N146), 
        .C1(N502), .Y(N497) );
  NOR2X2TF U218 ( .A(N338), .B(N955), .Y(N350) );
  NOR2X2TF U219 ( .A(N347), .B(N969), .Y(N383) );
  NOR3X2TF U220 ( .A(N110), .B(N604), .C(N631), .Y(N617) );
  INVX2TF U221 ( .A(N505), .Y(N126) );
  INVX2TF U222 ( .A(N505), .Y(N127) );
  INVX2TF U223 ( .A(N799), .Y(N130) );
  INVX2TF U224 ( .A(N799), .Y(N131) );
  NAND2X2TF U225 ( .A(N123), .B(N761), .Y(N454) );
  AOI21X2TF U226 ( .A0(N940), .A1(N920), .B0(N217), .Y(N934) );
  AOI211XLTF U227 ( .A0(N825), .A1(N824), .B0(OPER_A[2]), .C0(N915), .Y(N826)
         );
  OAI32XLTF U228 ( .A0(OPER_A[8]), .A1(N897), .A2(N915), .B0(N896), .B1(N895), 
        .Y(N898) );
  OAI32XLTF U229 ( .A0(OPER_A[10]), .A1(N916), .A2(N915), .B0(N914), .B1(N913), 
        .Y(N917) );
  OAI32XLTF U230 ( .A0(OPER_A[6]), .A1(N875), .A2(N915), .B0(N874), .B1(N873), 
        .Y(N876) );
  INVXLTF U231 ( .A(N915), .Y(N912) );
  INVX2TF U232 ( .A(DP_OP_333_124_4748_N57), .Y(N132) );
  CLKBUFX2TF U233 ( .A(N190), .Y(N133) );
  CLKBUFX2TF U234 ( .A(N257), .Y(N190) );
  NOR3XLTF U235 ( .A(N73), .B(N909), .C(N970), .Y(N819) );
  NAND2X2TF U236 ( .A(N968), .B(N928), .Y(N909) );
  AOI21XLTF U237 ( .A0(N820), .A1(N374), .B0(N373), .Y(N376) );
  AOI21XLTF U238 ( .A0(N822), .A1(N821), .B0(N820), .Y(N828) );
  INVXLTF U239 ( .A(N820), .Y(N377) );
  NOR3BX4TF U240 ( .AN(N385), .B(N382), .C(N125), .Y(N513) );
  AOI222X4TF U241 ( .A0(XTEMP[9]), .A1(X_IN[9]), .B0(XTEMP[9]), .B1(N478), 
        .C0(X_IN[9]), .C1(N478), .Y(N487) );
  AOI222X4TF U242 ( .A0(N175), .A1(N488), .B0(N175), .B1(N464), .C0(N488), 
        .C1(N464), .Y(N478) );
  OAI31XLTF U243 ( .A0(OPER_A[1]), .A1(N915), .A2(OPER_A[0]), .B0(N830), .Y(
        N831) );
  OAI21X2TF U244 ( .A0(N142), .A1(N107), .B0(N243), .Y(OPER_A[1]) );
  INVX2TF U245 ( .A(N123), .Y(N134) );
  NAND2X2TF U246 ( .A(N761), .B(N134), .Y(N558) );
  NOR2X4TF U247 ( .A(N386), .B(N767), .Y(N805) );
  AOI22XLTF U248 ( .A0(DIVISION_HEAD[5]), .A1(N87), .B0(X_IN[7]), .B1(N805), 
        .Y(N388) );
  AOI22XLTF U249 ( .A0(X_IN[10]), .A1(N130), .B0(X_IN[11]), .B1(N805), .Y(N427) );
  NOR4X2TF U250 ( .A(N647), .B(N942), .C(N366), .D(N365), .Y(N641) );
  NOR2X2TF U251 ( .A(N338), .B(N603), .Y(N565) );
  NOR2BX2TF U252 ( .AN(N543), .B(N383), .Y(N628) );
  INVX2TF U253 ( .A(N135), .Y(N136) );
  INVX2TF U254 ( .A(N135), .Y(N137) );
  AOI22X2TF U255 ( .A0(N345), .A1(N343), .B0(N939), .B1(N346), .Y(N921) );
  CLKBUFX2TF U256 ( .A(N1011), .Y(N138) );
  NOR2X1TF U257 ( .A(N115), .B(N189), .Y(N1011) );
  XNOR2X1TF U258 ( .A(OPER_A[12]), .B(ADD_X_132_1_N2), .Y(N139) );
  CMPR32X2TF U259 ( .A(OPER_A[7]), .B(OPER_B[7]), .C(ADD_X_132_1_N7), .CO(
        ADD_X_132_1_N6), .S(SUM_AB[7]) );
  CMPR32X2TF U260 ( .A(OPER_A[6]), .B(OPER_B[6]), .C(ADD_X_132_1_N8), .CO(
        ADD_X_132_1_N7), .S(SUM_AB[6]) );
  XNOR2X2TF U261 ( .A(N139), .B(OPER_B[12]), .Y(SUM_AB[12]) );
  AOI222XLTF U262 ( .A0(DIVISION_HEAD[1]), .A1(DIVISION_HEAD[0]), .B0(
        DIVISION_HEAD[1]), .B1(N314), .C0(DIVISION_HEAD[0]), .C1(N313), .Y(
        N316) );
  AOI32X1TF U263 ( .A0(N119), .A1(N56), .A2(N563), .B0(N617), .B1(N73), .Y(
        N544) );
  AOI22X1TF U264 ( .A0(N73), .A1(N162), .B0(POST_WORK), .B1(N109), .Y(N241) );
  NAND2X1TF U265 ( .A(N313), .B(N655), .Y(N315) );
  OAI31X1TF U266 ( .A0(N969), .A1(N948), .A2(N947), .B0(N946), .Y(N949) );
  NAND2X1TF U267 ( .A(N477), .B(N476), .Y(N486) );
  NOR2X1TF U268 ( .A(SUM_AB[8]), .B(N462), .Y(N477) );
  NOR2X1TF U269 ( .A(SUM_AB[10]), .B(N486), .Y(N499) );
  OA22X1TF U270 ( .A0(N767), .A1(N557), .B0(N762), .B1(N763), .Y(N305) );
  INVX2TF U271 ( .A(N928), .Y(N217) );
  OAI21X1TF U272 ( .A0(N947), .A1(N609), .B0(N646), .Y(N960) );
  NAND2X1TF U273 ( .A(Y_IN[1]), .B(Y_IN[0]), .Y(N314) );
  NAND2X1TF U274 ( .A(N564), .B(N346), .Y(N915) );
  NOR2X2TF U275 ( .A(N217), .B(N110), .Y(N903) );
  OR2X2TF U276 ( .A(N960), .B(N197), .Y(N928) );
  NOR2X1TF U277 ( .A(\INDEX[2] ), .B(N620), .Y(N308) );
  NAND2X1TF U278 ( .A(N129), .B(N128), .Y(N620) );
  OAI21X1TF U279 ( .A0(DIVISION_HEAD[12]), .A1(N548), .B0(N337), .Y(N947) );
  AOI2BB1X1TF U280 ( .A0N(DIVISION_HEAD[6]), .A1N(N326), .B0(Y_IN[6]), .Y(N324) );
  AOI2BB1X1TF U281 ( .A0N(DIVISION_HEAD[4]), .A1N(N322), .B0(Y_IN[4]), .Y(N320) );
  NAND2X1TF U282 ( .A(PRE_WORK), .B(N120), .Y(N386) );
  AOI211X1TF U283 ( .A0(Y_IN[11]), .A1(N301), .B0(Y_IN[12]), .C0(N282), .Y(
        N765) );
  CLKBUFX2TF U284 ( .A(N969), .Y(N189) );
  NAND2X1TF U285 ( .A(N911), .B(N903), .Y(N931) );
  AOI2BB1X1TF U286 ( .A0N(N607), .A1N(N342), .B0(N961), .Y(N197) );
  NOR2X1TF U287 ( .A(PRE_WORK), .B(N339), .Y(N341) );
  NAND2X1TF U288 ( .A(N122), .B(N148), .Y(N604) );
  NOR2X1TF U289 ( .A(N124), .B(N627), .Y(N339) );
  CLKBUFX2TF U290 ( .A(Y_IN[5]), .Y(N192) );
  NAND2X1TF U291 ( .A(N140), .B(N149), .Y(N338) );
  NAND2X1TF U292 ( .A(N454), .B(N460), .Y(N471) );
  NAND2X2TF U293 ( .A(N546), .B(N385), .Y(N460) );
  CLKBUFX2TF U294 ( .A(N780), .Y(N191) );
  NAND2X1TF U295 ( .A(N121), .B(N122), .Y(N955) );
  AND2X2TF U296 ( .A(ALU_START), .B(N133), .Y(N218) );
  NAND2X1TF U297 ( .A(N565), .B(N383), .Y(N609) );
  NAND2X2TF U298 ( .A(N219), .B(ALU_START), .Y(N969) );
  NAND2X1TF U299 ( .A(N174), .B(N364), .Y(N347) );
  NAND2X1TF U300 ( .A(N124), .B(N308), .Y(N364) );
  NAND2X1TF U301 ( .A(N121), .B(N163), .Y(N603) );
  AND2X2TF U302 ( .A(N196), .B(ALU_TYPE[1]), .Y(N219) );
  AOI211X1TF U303 ( .A0(N218), .A1(N607), .B0(N944), .C0(N606), .Y(N610) );
  NOR3X1TF U304 ( .A(N605), .B(N604), .C(N775), .Y(N606) );
  OR3X1TF U305 ( .A(N881), .B(N880), .C(N212), .Y(N676) );
  OAI2BB2XLTF U306 ( .B0(N882), .B1(N970), .A0N(C152_DATA4_6), .A1N(N104), .Y(
        N212) );
  OAI2BB2XLTF U307 ( .B0(N879), .B1(N923), .A0N(N217), .A1N(OPER_B[6]), .Y(
        N880) );
  INVX2TF U308 ( .A(N460), .Y(N475) );
  AOI32X1TF U309 ( .A0(N968), .A1(N114), .A2(N967), .B0(N119), .B1(N114), .Y(
        N1018) );
  NOR2BX2TF U310 ( .AN(N546), .B(N556), .Y(N812) );
  NOR2X1TF U311 ( .A(N174), .B(N599), .Y(N352) );
  NAND2X1TF U312 ( .A(N959), .B(DP_OP_333_124_4748_N57), .Y(N649) );
  INVX2TF U313 ( .A(N363), .Y(N761) );
  NAND2X1TF U314 ( .A(N383), .B(N959), .Y(N363) );
  NAND2X1TF U315 ( .A(N903), .B(N870), .Y(N893) );
  NOR2X1TF U316 ( .A(N56), .B(N909), .Y(N905) );
  AND2X2TF U317 ( .A(N218), .B(PRE_WORK), .Y(DP_OP_333_124_4748_N57) );
  AOI21X1TF U318 ( .A0(N948), .A1(N966), .B0(N362), .Y(N968) );
  NAND2X1TF U319 ( .A(N140), .B(STEP[3]), .Y(N631) );
  NOR2X2TF U320 ( .A(N338), .B(N604), .Y(N959) );
  NAND2X1TF U321 ( .A(N339), .B(N174), .Y(N344) );
  NAND3X1TF U322 ( .A(N961), .B(N969), .C(N599), .Y(N646) );
  INVX2TF U323 ( .A(N218), .Y(N961) );
  NOR3BX1TF U324 ( .AN(ALU_TYPE[0]), .B(ALU_TYPE[1]), .C(ALU_TYPE[2]), .Y(N257) );
  AO22X1TF U325 ( .A0(N371), .A1(XTEMP[12]), .B0(N359), .B1(N964), .Y(N722) );
  AOI32X1TF U326 ( .A0(N966), .A1(N360), .A2(N957), .B0(N972), .B1(N360), .Y(
        N361) );
  NAND2X1TF U327 ( .A(N945), .B(DP_OP_333_124_4748_N57), .Y(N634) );
  NAND2X1TF U328 ( .A(N642), .B(N113), .Y(N614) );
  NAND2X1TF U329 ( .A(N104), .B(C152_DATA4_8), .Y(N213) );
  AOI32X1TF U330 ( .A0(N117), .A1(DIVISION_HEAD[4]), .A2(N748), .B0(N471), 
        .B1(DIVISION_HEAD[4]), .Y(N392) );
  OAI22X1TF U331 ( .A0(N528), .A1(N93), .B0(N488), .B1(N95), .Y(N489) );
  INVX2TF U332 ( .A(N1014), .Y(N1009) );
  OAI2BB2XLTF U333 ( .B0(N56), .B1(N970), .A0N(N970), .A1N(N56), .Y(N973) );
  NAND2X1TF U334 ( .A(N646), .B(N94), .Y(N943) );
  NAND2X1TF U335 ( .A(N565), .B(DP_OP_333_124_4748_N57), .Y(N394) );
  INVX2TF U336 ( .A(N112), .Y(N775) );
  NOR2X2TF U337 ( .A(N761), .B(N191), .Y(N759) );
  NAND2X1TF U338 ( .A(N350), .B(N112), .Y(N543) );
  NOR2X1TF U339 ( .A(N955), .B(N631), .Y(N563) );
  OAI21X2TF U340 ( .A0(N151), .A1(N107), .B0(N242), .Y(OPER_A[0]) );
  NOR2X1TF U341 ( .A(N604), .B(N953), .Y(N564) );
  NAND2X1TF U342 ( .A(STEP[2]), .B(N149), .Y(N953) );
  OAI32X1TF U343 ( .A0(N648), .A1(N177), .A2(N943), .B0(N147), .B1(N649), .Y(
        N694) );
  OAI21X1TF U344 ( .A0(N174), .A1(N647), .B0(N646), .Y(N695) );
  AOI22X1TF U345 ( .A0(N542), .A1(N73), .B0(N541), .B1(N540), .Y(N707) );
  INVX2TF U346 ( .A(N542), .Y(N540) );
  OAI31X1TF U347 ( .A0(N539), .A1(N538), .A2(N537), .B0(N536), .Y(N541) );
  AOI211X1TF U348 ( .A0(N535), .A1(XTEMP[12]), .B0(N534), .C0(N533), .Y(N536)
         );
  OAI31X1TF U349 ( .A0(DIVISION_HEAD[1]), .A1(N532), .A2(N146), .B0(N531), .Y(
        N535) );
  AOI22X1TF U350 ( .A0(N530), .A1(N529), .B0(XTEMP[11]), .B1(N161), .Y(N531)
         );
  OAI22X1TF U351 ( .A0(DIVISION_HEAD[0]), .A1(N528), .B0(DIVISION_REMA[8]), 
        .B1(N175), .Y(N529) );
  INVX2TF U352 ( .A(N538), .Y(N530) );
  NOR2X1TF U353 ( .A(XTEMP[11]), .B(N161), .Y(N532) );
  OAI22X1TF U354 ( .A0(DIVISION_HEAD[12]), .A1(N145), .B0(XTEMP[12]), .B1(N147), .Y(N537) );
  OAI21X1TF U355 ( .A0(XTEMP[11]), .A1(N161), .B0(N527), .Y(N538) );
  AOI22X1TF U356 ( .A0(DIVISION_HEAD[0]), .A1(N528), .B0(DIVISION_HEAD[1]), 
        .B1(N146), .Y(N527) );
  AOI21X1TF U357 ( .A0(DIVISION_HEAD[11]), .A1(N166), .B0(N526), .Y(N539) );
  AOI211X1TF U358 ( .A0(DIVISION_REMA[6]), .A1(N153), .B0(N525), .C0(N524), 
        .Y(N526) );
  NOR2X1TF U359 ( .A(DIVISION_HEAD[11]), .B(N166), .Y(N524) );
  AOI21X1TF U360 ( .A0(DIVISION_HEAD[9]), .A1(N165), .B0(N522), .Y(N523) );
  AOI211X1TF U361 ( .A0(DIVISION_REMA[4]), .A1(N152), .B0(N521), .C0(N520), 
        .Y(N522) );
  NOR2X1TF U362 ( .A(DIVISION_HEAD[9]), .B(N165), .Y(N520) );
  AOI21X1TF U363 ( .A0(DIVISION_HEAD[7]), .A1(N164), .B0(N518), .Y(N519) );
  AOI211X1TF U364 ( .A0(N517), .A1(DIVISION_REMA[2]), .B0(N516), .C0(N515), 
        .Y(N518) );
  NOR2X1TF U365 ( .A(DIVISION_HEAD[7]), .B(N164), .Y(N516) );
  OAI21X1TF U366 ( .A0(DIVISION_HEAD[5]), .A1(N158), .B0(N514), .Y(N517) );
  OAI211X1TF U367 ( .A0(DIVISION_REMA[1]), .A1(N142), .B0(DIVISION_REMA[0]), 
        .C0(N151), .Y(N514) );
  OAI21X1TF U368 ( .A0(N380), .A1(N162), .B0(N379), .Y(N720) );
  OAI22X1TF U369 ( .A0(N111), .A1(N377), .B0(N762), .B1(N639), .Y(N378) );
  OAI211X1TF U370 ( .A0(N372), .A1(N821), .B0(N611), .C0(N639), .Y(N373) );
  OAI21X1TF U371 ( .A0(N949), .A1(N968), .B0(N951), .Y(N950) );
  OR4X2TF U372 ( .A(N944), .B(N943), .C(N942), .D(N941), .Y(N951) );
  OAI22X1TF U373 ( .A0(N111), .A1(N939), .B0(N938), .B1(N972), .Y(N941) );
  OAI21X1TF U374 ( .A0(N596), .A1(N585), .B0(N584), .Y(N702) );
  AOI31X1TF U375 ( .A0(N583), .A1(N588), .A2(N590), .B0(N582), .Y(N585) );
  OAI22X1TF U376 ( .A0(N128), .A1(N581), .B0(N592), .B1(N588), .Y(N582) );
  OAI21X1TF U377 ( .A0(N128), .A1(N619), .B0(N618), .Y(N699) );
  AOI31X1TF U378 ( .A0(N617), .A1(N620), .A2(N616), .B0(N615), .Y(N618) );
  OAI32X1TF U379 ( .A0(N628), .A1(N629), .A2(N620), .B0(N616), .B1(N628), .Y(
        N615) );
  AOI22X1TF U380 ( .A0(N596), .A1(N92), .B0(N580), .B1(N579), .Y(N703) );
  AOI211X1TF U381 ( .A0(N594), .A1(N156), .B0(N578), .C0(N789), .Y(N580) );
  AOI21X1TF U382 ( .A0(N577), .A1(N775), .B0(N179), .Y(N578) );
  OAI21X1TF U383 ( .A0(N129), .A1(N619), .B0(N307), .Y(N726) );
  OAI21X1TF U384 ( .A0(N306), .A1(N382), .B0(N619), .Y(N307) );
  AOI32X1TF U385 ( .A0(N628), .A1(N634), .A2(N375), .B0(N156), .B1(N634), .Y(
        N306) );
  OAI31X1TF U386 ( .A0(N629), .A1(N628), .A2(N627), .B0(N626), .Y(N698) );
  AOI22X1TF U387 ( .A0(\INDEX[2] ), .A1(N625), .B0(N624), .B1(N623), .Y(N626)
         );
  OAI21X1TF U388 ( .A0(N622), .A1(N628), .B0(N621), .Y(N625) );
  AOI32X1TF U389 ( .A0(N310), .A1(N124), .A2(N617), .B0(N185), .B1(N309), .Y(
        N312) );
  NOR2X1TF U390 ( .A(N629), .B(N623), .Y(N621) );
  AOI21X1TF U391 ( .A0(\INDEX[2] ), .A1(N624), .B0(N375), .Y(N623) );
  INVX2TF U392 ( .A(N619), .Y(N629) );
  INVX2TF U393 ( .A(N616), .Y(N624) );
  OAI211X1TF U394 ( .A0(N111), .A1(N368), .B0(N644), .C0(N367), .Y(N721) );
  AOI22X1TF U395 ( .A0(STEP[3]), .A1(N641), .B0(N374), .B1(N573), .Y(N367) );
  OAI211X1TF U396 ( .A0(N178), .A1(N614), .B0(N630), .C0(N613), .Y(N700) );
  AOI21X1TF U397 ( .A0(N641), .A1(N148), .B0(N612), .Y(N613) );
  NOR3X1TF U398 ( .A(STEP[3]), .B(N111), .C(N603), .Y(N944) );
  AOI211X1TF U399 ( .A0(N822), .A1(N374), .B0(N371), .C0(N370), .Y(N611) );
  AOI21X1TF U400 ( .A0(N384), .A1(N369), .B0(N775), .Y(N370) );
  NOR2X1TF U401 ( .A(N110), .B(N821), .Y(N374) );
  OAI22X1TF U402 ( .A0(N90), .A1(N597), .B0(N596), .B1(N595), .Y(N701) );
  AOI21X1TF U403 ( .A0(\INDEX[2] ), .A1(N594), .B0(N593), .Y(N595) );
  OAI22X1TF U404 ( .A0(N592), .A1(N591), .B0(N590), .B1(N589), .Y(N593) );
  INVX2TF U405 ( .A(N587), .Y(N592) );
  AOI21X1TF U406 ( .A0(N588), .A1(N587), .B0(N586), .Y(N597) );
  OAI211X1TF U407 ( .A0(N645), .A1(N140), .B0(N644), .C0(N643), .Y(N696) );
  NOR2X1TF U408 ( .A(N648), .B(N361), .Y(N644) );
  OAI21X1TF U409 ( .A0(N350), .A1(N259), .B0(N119), .Y(N360) );
  INVX2TF U410 ( .A(N649), .Y(N648) );
  OAI22X1TF U411 ( .A0(N163), .A1(N953), .B0(N821), .B1(N966), .Y(N637) );
  AOI211X1TF U412 ( .A0(N641), .A1(N163), .B0(N636), .C0(N635), .Y(N640) );
  INVX2TF U413 ( .A(N260), .Y(N633) );
  AOI31X1TF U414 ( .A0(N955), .A1(N369), .A2(N384), .B0(N775), .Y(N260) );
  AOI21X1TF U415 ( .A0(N120), .A1(N602), .B0(N601), .Y(N630) );
  OAI21X1TF U416 ( .A0(N600), .A1(N599), .B0(N598), .Y(N601) );
  OAI22X1TF U417 ( .A0(N596), .A1(N576), .B0(N575), .B1(N188), .Y(N704) );
  AOI21X1TF U418 ( .A0(N591), .A1(N587), .B0(N586), .Y(N575) );
  OAI21X1TF U419 ( .A0(N90), .A1(N590), .B0(N583), .Y(N589) );
  INVX2TF U420 ( .A(N614), .Y(N583) );
  INVX2TF U421 ( .A(N596), .Y(N579) );
  OAI31X1TF U422 ( .A0(N605), .A1(N604), .A2(N775), .B0(N577), .Y(N587) );
  OAI32X1TF U423 ( .A0(N574), .A1(N822), .A2(N573), .B0(N119), .B1(N574), .Y(
        N577) );
  INVX2TF U424 ( .A(N572), .Y(N574) );
  AOI21X1TF U425 ( .A0(N594), .A1(N185), .B0(N571), .Y(N576) );
  AOI32X1TF U426 ( .A0(N565), .A1(N113), .A2(N178), .B0(N959), .B1(N112), .Y(
        N567) );
  AOI31X1TF U427 ( .A0(N119), .A1(N822), .A2(N821), .B0(N943), .Y(N568) );
  INVX2TF U428 ( .A(N581), .Y(N594) );
  AOI22X1TF U429 ( .A0(N902), .A1(N903), .B0(N217), .B1(OPER_B[8]), .Y(N214)
         );
  OAI21X1TF U430 ( .A0(N901), .A1(N159), .B0(N900), .Y(N902) );
  AOI211X1TF U431 ( .A0(N919), .A1(OPER_B[9]), .B0(N899), .C0(N898), .Y(N900)
         );
  AOI21X1TF U432 ( .A0(N912), .A1(N897), .B0(N911), .Y(N895) );
  NOR3X1TF U433 ( .A(N910), .B(OPER_B[8]), .C(N894), .Y(N899) );
  AOI21X1TF U434 ( .A0(N894), .A1(N921), .B0(N920), .Y(N901) );
  OAI211X1TF U435 ( .A0(N1009), .A1(N996), .B0(N995), .C0(N994), .Y(N662) );
  AOI22X1TF U436 ( .A0(DIVISION_HEAD[7]), .A1(N1011), .B0(ZTEMP[7]), .B1(N116), 
        .Y(N995) );
  OAI211X1TF U437 ( .A0(N1009), .A1(N990), .B0(N989), .C0(N988), .Y(N664) );
  AOI22X1TF U438 ( .A0(DIVISION_HEAD[5]), .A1(N138), .B0(ZTEMP[5]), .B1(N116), 
        .Y(N989) );
  OAI211X1TF U439 ( .A0(N1009), .A1(N984), .B0(N983), .C0(N982), .Y(N666) );
  AOI22X1TF U440 ( .A0(DIVISION_HEAD[3]), .A1(N138), .B0(ZTEMP[3]), .B1(N116), 
        .Y(N983) );
  AOI22X1TF U441 ( .A0(SUM_AB[2]), .A1(N81), .B0(N979), .B1(N1014), .Y(N980)
         );
  AOI22X1TF U442 ( .A0(DIVISION_HEAD[2]), .A1(N138), .B0(ZTEMP[2]), .B1(N115), 
        .Y(N981) );
  AOI22X1TF U443 ( .A0(SUM_AB[6]), .A1(N81), .B0(N991), .B1(N1014), .Y(N992)
         );
  AOI22X1TF U444 ( .A0(DIVISION_HEAD[6]), .A1(N138), .B0(ZTEMP[6]), .B1(N116), 
        .Y(N993) );
  AOI22X1TF U445 ( .A0(SUM_AB[4]), .A1(N81), .B0(N985), .B1(N1014), .Y(N986)
         );
  AOI22X1TF U446 ( .A0(DIVISION_HEAD[4]), .A1(N138), .B0(ZTEMP[4]), .B1(N115), 
        .Y(N987) );
  AOI22X1TF U447 ( .A0(SUM_AB[1]), .A1(N81), .B0(N976), .B1(N1014), .Y(N977)
         );
  AOI22X1TF U448 ( .A0(DIVISION_HEAD[1]), .A1(N138), .B0(ZTEMP[1]), .B1(N116), 
        .Y(N978) );
  OAI21X1TF U449 ( .A0(N450), .A1(N449), .B0(N460), .Y(N451) );
  AOI22X1TF U450 ( .A0(DIVISION_HEAD[11]), .A1(N88), .B0(X_IN[12]), .B1(N131), 
        .Y(N445) );
  AOI22X1TF U451 ( .A0(SUM_AB[6]), .A1(N126), .B0(N493), .B1(N991), .Y(N447)
         );
  OAI22X1TF U452 ( .A0(N144), .A1(N93), .B0(N442), .B1(N95), .Y(N450) );
  AOI22X1TF U453 ( .A0(SUM_AB[8]), .A1(N81), .B0(N997), .B1(N1014), .Y(N998)
         );
  AOI22X1TF U454 ( .A0(DIVISION_HEAD[8]), .A1(N138), .B0(ZTEMP[8]), .B1(N115), 
        .Y(N999) );
  OAI211X1TF U455 ( .A0(N1009), .A1(N1002), .B0(N1001), .C0(N1000), .Y(N660)
         );
  AOI22X1TF U456 ( .A0(DIVISION_HEAD[9]), .A1(N1011), .B0(ZTEMP[9]), .B1(N116), 
        .Y(N1001) );
  INVX2TF U457 ( .A(N881), .Y(N209) );
  AOI31X1TF U458 ( .A0(N835), .A1(N834), .A2(N833), .B0(N923), .Y(N837) );
  AOI32X1TF U459 ( .A0(N832), .A1(OPER_B[2]), .A2(N921), .B0(N920), .B1(
        OPER_B[2]), .Y(N833) );
  AOI22X1TF U460 ( .A0(N919), .A1(OPER_B[3]), .B0(OPER_A[2]), .B1(N831), .Y(
        N834) );
  AOI31X1TF U461 ( .A0(N921), .A1(N155), .A2(N827), .B0(N826), .Y(N835) );
  AOI211X1TF U462 ( .A0(N217), .A1(OPER_B[10]), .B0(N926), .C0(N927), .Y(N215)
         );
  AOI21X1TF U463 ( .A0(N974), .A1(N970), .B0(N909), .Y(N927) );
  AOI21X1TF U464 ( .A0(N925), .A1(N924), .B0(N923), .Y(N926) );
  AOI32X1TF U465 ( .A0(N922), .A1(OPER_B[10]), .A2(N921), .B0(N920), .B1(
        OPER_B[10]), .Y(N924) );
  AOI211X1TF U466 ( .A0(N919), .A1(OPER_B[11]), .B0(N918), .C0(N917), .Y(N925)
         );
  AOI21X1TF U467 ( .A0(N912), .A1(N916), .B0(N911), .Y(N913) );
  NOR3X1TF U468 ( .A(N910), .B(OPER_B[10]), .C(N922), .Y(N918) );
  OAI22X1TF U469 ( .A0(N475), .A1(N474), .B0(N473), .B1(N175), .Y(N711) );
  AOI211X1TF U470 ( .A0(N997), .A1(N493), .B0(N470), .C0(N469), .Y(N474) );
  OAI211X1TF U471 ( .A0(N468), .A1(N608), .B0(N467), .C0(N466), .Y(N469) );
  AOI22X1TF U472 ( .A0(XTEMP[9]), .A1(N88), .B0(N798), .B1(SUM_AB[12]), .Y(
        N466) );
  NOR2X1TF U473 ( .A(DIVISION_HEAD[12]), .B(N472), .Y(N465) );
  AOI22X1TF U474 ( .A0(X_IN[8]), .A1(N464), .B0(INTADD_0_N1), .B1(N488), .Y(
        N472) );
  OAI22X1TF U475 ( .A0(N141), .A1(N93), .B0(N463), .B1(N95), .Y(N470) );
  AOI211X1TF U476 ( .A0(OPER_B[6]), .A1(N878), .B0(N877), .C0(N876), .Y(N879)
         );
  AOI21X1TF U477 ( .A0(N912), .A1(N875), .B0(N911), .Y(N873) );
  OAI31X1TF U478 ( .A0(N910), .A1(OPER_B[6]), .A2(N872), .B0(N871), .Y(N877)
         );
  AOI21X1TF U479 ( .A0(OPER_B[7]), .A1(N870), .B0(N869), .Y(N871) );
  OAI21X1TF U480 ( .A0(N910), .A1(N868), .B0(N867), .Y(N878) );
  AOI32X1TF U481 ( .A0(N431), .A1(N460), .A2(N430), .B0(N475), .B1(N152), .Y(
        N715) );
  AOI211X1TF U482 ( .A0(N493), .A1(N985), .B0(N429), .C0(N428), .Y(N430) );
  AOI22X1TF U483 ( .A0(DIVISION_HEAD[9]), .A1(N87), .B0(X_IN[9]), .B1(N99), 
        .Y(N426) );
  OAI22X1TF U484 ( .A0(N143), .A1(N93), .B0(N152), .B1(N454), .Y(N429) );
  AOI32X1TF U485 ( .A0(N393), .A1(N392), .A2(N391), .B0(N475), .B1(N392), .Y(
        N719) );
  OAI211X1TF U486 ( .A0(N389), .A1(N558), .B0(N388), .C0(N387), .Y(N390) );
  AOI22X1TF U487 ( .A0(X_IN[6]), .A1(N131), .B0(X_IN[5]), .B1(N99), .Y(N387)
         );
  AOI22X1TF U488 ( .A0(DIVISION_HEAD[3]), .A1(N734), .B0(SUM_AB[0]), .B1(N381), 
        .Y(N393) );
  AOI32X1TF U489 ( .A0(N412), .A1(N460), .A2(N411), .B0(N475), .B1(N150), .Y(
        N717) );
  AOI211X1TF U490 ( .A0(DIVISION_HEAD[7]), .A1(N88), .B0(N410), .C0(N409), .Y(
        N411) );
  OAI211X1TF U491 ( .A0(N95), .A1(N748), .B0(N408), .C0(N407), .Y(N409) );
  AOI21X1TF U492 ( .A0(N493), .A1(N979), .B0(N406), .Y(N407) );
  OAI22X1TF U493 ( .A0(N142), .A1(N89), .B0(N150), .B1(N454), .Y(N406) );
  AOI22X1TF U494 ( .A0(X_IN[1]), .A1(N444), .B0(N798), .B1(SUM_AB[6]), .Y(N408) );
  OAI21X1TF U495 ( .A0(N500), .A1(N747), .B0(N403), .Y(N410) );
  AOI22X1TF U496 ( .A0(X_IN[8]), .A1(N131), .B0(X_IN[7]), .B1(N99), .Y(N403)
         );
  AOI32X1TF U497 ( .A0(N402), .A1(N460), .A2(N401), .B0(N475), .B1(N142), .Y(
        N718) );
  AOI211X1TF U498 ( .A0(N493), .A1(N976), .B0(N400), .C0(N399), .Y(N401) );
  OAI211X1TF U499 ( .A0(N558), .A1(N432), .B0(N398), .C0(N397), .Y(N399) );
  AOI21X1TF U500 ( .A0(DIVISION_HEAD[4]), .A1(N734), .B0(N396), .Y(N397) );
  OAI22X1TF U501 ( .A0(N142), .A1(N454), .B0(N748), .B1(N608), .Y(N396) );
  AOI22X1TF U502 ( .A0(DIVISION_HEAD[6]), .A1(N88), .B0(X_IN[7]), .B1(N130), 
        .Y(N398) );
  OAI22X1TF U503 ( .A0(N463), .A1(N395), .B0(N488), .B1(N747), .Y(N400) );
  OAI22X1TF U504 ( .A0(N513), .A1(N485), .B0(N484), .B1(N528), .Y(N710) );
  AOI211X1TF U505 ( .A0(SUM_AB[9]), .A1(N127), .B0(N482), .C0(N481), .Y(N485)
         );
  OAI211X1TF U506 ( .A0(N1002), .A1(N507), .B0(N480), .C0(N479), .Y(N481) );
  AOI22X1TF U507 ( .A0(XTEMP[10]), .A1(N88), .B0(X_IN[7]), .B1(N800), .Y(N480)
         );
  OAI22X1TF U508 ( .A0(N175), .A1(N93), .B0(N488), .B1(N608), .Y(N482) );
  AOI32X1TF U509 ( .A0(N461), .A1(N460), .A2(N459), .B0(N475), .B1(N141), .Y(
        N712) );
  OAI211X1TF U510 ( .A0(N507), .A1(N996), .B0(N456), .C0(N455), .Y(N457) );
  AOI22X1TF U511 ( .A0(DIVISION_HEAD[12]), .A1(N87), .B0(X_IN[12]), .B1(N98), 
        .Y(N455) );
  AOI22X1TF U512 ( .A0(DIVISION_HEAD[11]), .A1(N804), .B0(DIVISION_HEAD[10]), 
        .B1(N125), .Y(N456) );
  OAI22X1TF U513 ( .A0(N463), .A1(N608), .B0(N558), .B1(N498), .Y(N458) );
  AOI22X1TF U514 ( .A0(SUM_AB[10]), .A1(N82), .B0(N1003), .B1(N1014), .Y(N1004) );
  AOI22X1TF U515 ( .A0(DIVISION_HEAD[10]), .A1(N138), .B0(ZTEMP[10]), .B1(N116), .Y(N1005) );
  AOI32X1TF U516 ( .A0(N797), .A1(N814), .A2(N796), .B0(N812), .B1(N172), .Y(
        N684) );
  AOI21X1TF U517 ( .A0(N795), .A1(N1003), .B0(N794), .Y(N796) );
  AOI22X1TF U518 ( .A0(X_IN[2]), .A1(N99), .B0(X_IN[4]), .B1(N805), .Y(N790)
         );
  AOI22X1TF U519 ( .A0(DIVISION_HEAD[0]), .A1(N125), .B0(DIVISION_HEAD[1]), 
        .B1(N804), .Y(N791) );
  AOI22X1TF U520 ( .A0(Y_IN[10]), .A1(N789), .B0(X_IN[3]), .B1(N131), .Y(N792)
         );
  AOI22X1TF U521 ( .A0(N798), .A1(SUM_AB[1]), .B0(SUM_AB[10]), .B1(N137), .Y(
        N797) );
  OAI22X1TF U522 ( .A0(N513), .A1(N496), .B0(N495), .B1(N146), .Y(N709) );
  AOI21X1TF U523 ( .A0(N493), .A1(N1003), .B0(N492), .Y(N496) );
  OAI211X1TF U524 ( .A0(N500), .A1(N608), .B0(N491), .C0(N490), .Y(N492) );
  AOI22X1TF U525 ( .A0(XTEMP[11]), .A1(N88), .B0(SUM_AB[10]), .B1(N126), .Y(
        N491) );
  AOI21X1TF U526 ( .A0(SUM_AB[10]), .A1(N486), .B0(N499), .Y(N1003) );
  AOI22X1TF U527 ( .A0(N191), .A1(N145), .B0(N779), .B1(N778), .Y(N686) );
  AOI211X1TF U528 ( .A0(DIVISION_REMA[7]), .A1(N734), .B0(N777), .C0(N776), 
        .Y(N779) );
  OAI211X1TF U529 ( .A0(N167), .A1(N775), .B0(N774), .C0(N773), .Y(N776) );
  AOI22X1TF U530 ( .A0(N772), .A1(N771), .B0(N997), .B1(N795), .Y(N773) );
  AOI21X1TF U531 ( .A0(SUM_AB[8]), .A1(N462), .B0(N477), .Y(N997) );
  AOI32X1TF U532 ( .A0(N770), .A1(N769), .A2(N768), .B0(N767), .B1(N769), .Y(
        N771) );
  OAI32X1TF U533 ( .A0(N766), .A1(N765), .A2(X_IN[0]), .B0(N764), .B1(N766), 
        .Y(N769) );
  AOI22X1TF U534 ( .A0(DIVISION_REMA[8]), .A1(N761), .B0(SUM_AB[8]), .B1(N136), 
        .Y(N774) );
  AOI22X1TF U535 ( .A0(N475), .A1(N144), .B0(N441), .B1(N460), .Y(N714) );
  AOI21X1TF U536 ( .A0(DIVISION_HEAD[8]), .A1(N125), .B0(N434), .Y(N435) );
  OAI22X1TF U537 ( .A0(N144), .A1(N454), .B0(N507), .B1(N990), .Y(N434) );
  AOI22X1TF U538 ( .A0(DIVISION_HEAD[10]), .A1(N87), .B0(X_IN[10]), .B1(N98), 
        .Y(N437) );
  OAI22X1TF U539 ( .A0(N442), .A1(N608), .B0(N558), .B1(N476), .Y(N440) );
  OAI211X1TF U540 ( .A0(N1009), .A1(N1008), .B0(N1007), .C0(N1006), .Y(N658)
         );
  AOI22X1TF U541 ( .A0(DIVISION_HEAD[11]), .A1(N138), .B0(ZTEMP[11]), .B1(N116), .Y(N1007) );
  AOI32X1TF U542 ( .A0(N422), .A1(N460), .A2(N421), .B0(N475), .B1(N143), .Y(
        N716) );
  AOI211X1TF U543 ( .A0(DIVISION_HEAD[8]), .A1(N88), .B0(N420), .C0(N419), .Y(
        N421) );
  OAI211X1TF U544 ( .A0(N558), .A1(N452), .B0(N418), .C0(N417), .Y(N419) );
  AOI21X1TF U545 ( .A0(DIVISION_HEAD[6]), .A1(N734), .B0(N416), .Y(N417) );
  OAI22X1TF U546 ( .A0(N143), .A1(N454), .B0(N507), .B1(N984), .Y(N416) );
  OAI21X1TF U547 ( .A0(N502), .A1(N747), .B0(N413), .Y(N420) );
  AOI22X1TF U548 ( .A0(X_IN[8]), .A1(N99), .B0(X_IN[9]), .B1(N131), .Y(N413)
         );
  OAI21X1TF U549 ( .A0(N759), .A1(N178), .B0(N562), .Y(N705) );
  OAI22X1TF U550 ( .A0(N561), .A1(N560), .B0(N761), .B1(N778), .Y(N562) );
  AOI22X1TF U551 ( .A0(Y_IN[0]), .A1(N789), .B0(DIVISION_REMA[1]), .B1(N112), 
        .Y(N559) );
  AOI21X1TF U552 ( .A0(N111), .A1(N649), .B0(N975), .Y(N561) );
  INVX2TF U553 ( .A(SUM_AB[0]), .Y(N975) );
  OAI22X1TF U554 ( .A0(N191), .A1(N653), .B0(N759), .B1(N158), .Y(N693) );
  AOI21X1TF U555 ( .A0(SUM_AB[1]), .A1(N137), .B0(N652), .Y(N653) );
  AOI22X1TF U556 ( .A0(DIVISION_REMA[0]), .A1(N734), .B0(N795), .B1(N976), .Y(
        N650) );
  AOI21X1TF U557 ( .A0(SUM_AB[1]), .A1(SUM_AB[0]), .B0(N404), .Y(N976) );
  AOI22X1TF U558 ( .A0(Y_IN[1]), .A1(N789), .B0(DIVISION_REMA[2]), .B1(N113), 
        .Y(N651) );
  OAI22X1TF U559 ( .A0(N191), .A1(N739), .B0(N759), .B1(N168), .Y(N690) );
  AOI211X1TF U560 ( .A0(SUM_AB[4]), .A1(N137), .B0(N738), .C0(N737), .Y(N739)
         );
  OAI211X1TF U561 ( .A0(N736), .A1(N95), .B0(N755), .C0(N735), .Y(N737) );
  AOI22X1TF U562 ( .A0(DIVISION_REMA[5]), .A1(N113), .B0(N795), .B1(N985), .Y(
        N735) );
  AOI21X1TF U563 ( .A0(SUM_AB[4]), .A1(N423), .B0(N433), .Y(N985) );
  OAI22X1TF U564 ( .A0(N200), .A1(N802), .B0(N164), .B1(N93), .Y(N738) );
  OAI22X1TF U565 ( .A0(N191), .A1(N728), .B0(N759), .B1(N171), .Y(N692) );
  AOI211X1TF U566 ( .A0(SUM_AB[2]), .A1(N137), .B0(N727), .C0(N656), .Y(N728)
         );
  OAI211X1TF U567 ( .A0(N655), .A1(N95), .B0(N755), .C0(N654), .Y(N656) );
  AOI22X1TF U568 ( .A0(DIVISION_REMA[3]), .A1(N113), .B0(N795), .B1(N979), .Y(
        N654) );
  AOI21X1TF U569 ( .A0(SUM_AB[2]), .A1(N405), .B0(N415), .Y(N979) );
  NOR2X1TF U570 ( .A(SUM_AB[0]), .B(SUM_AB[1]), .Y(N404) );
  OAI22X1TF U571 ( .A0(N736), .A1(N802), .B0(N158), .B1(N93), .Y(N727) );
  OAI22X1TF U572 ( .A0(N191), .A1(N751), .B0(N759), .B1(N173), .Y(N688) );
  AOI211X1TF U573 ( .A0(N991), .A1(N795), .B0(N750), .C0(N749), .Y(N751) );
  OAI211X1TF U574 ( .A0(N748), .A1(N747), .B0(N755), .C0(N746), .Y(N749) );
  AOI22X1TF U575 ( .A0(DIVISION_REMA[7]), .A1(N112), .B0(SUM_AB[6]), .B1(N136), 
        .Y(N746) );
  INVX2TF U576 ( .A(N805), .Y(N747) );
  OAI21X1TF U577 ( .A0(N200), .A1(N95), .B0(N744), .Y(N750) );
  AOI22X1TF U578 ( .A0(Y_IN[6]), .A1(N789), .B0(DIVISION_REMA[5]), .B1(N734), 
        .Y(N744) );
  AOI21X1TF U579 ( .A0(SUM_AB[6]), .A1(N443), .B0(N453), .Y(N991) );
  INVX2TF U580 ( .A(N921), .Y(N910) );
  OAI211X1TF U581 ( .A0(N1018), .A1(N1017), .B0(N1016), .C0(N1015), .Y(N657)
         );
  AOI32X1TF U582 ( .A0(N1017), .A1(N1014), .A2(N1013), .B0(N1012), .B1(N1014), 
        .Y(N1015) );
  AOI211X4TF U583 ( .A0(N974), .A1(N973), .B0(N972), .C0(N115), .Y(N1014) );
  INVX2TF U584 ( .A(N968), .Y(N972) );
  AOI22X1TF U585 ( .A0(DIVISION_HEAD[12]), .A1(N138), .B0(ZTEMP[12]), .B1(N116), .Y(N1016) );
  OAI31X1TF U586 ( .A0(N966), .A1(N56), .A2(N970), .B0(N965), .Y(N967) );
  AOI31X1TF U587 ( .A0(N177), .A1(N56), .A2(N964), .B0(N963), .Y(N965) );
  AOI31X1TF U588 ( .A0(N959), .A1(N958), .A2(N957), .B0(N956), .Y(N962) );
  OAI31X1TF U589 ( .A0(N955), .A1(N954), .A2(N953), .B0(N952), .Y(N956) );
  OAI22X1TF U590 ( .A0(N513), .A1(N358), .B0(N357), .B1(N170), .Y(N723) );
  AOI211X1TF U591 ( .A0(N493), .A1(N1012), .B0(N355), .C0(N354), .Y(N358) );
  OAI31X1TF U592 ( .A0(XTEMP[12]), .A1(N356), .A2(N509), .B0(N353), .Y(N354)
         );
  INVX2TF U593 ( .A(N608), .Y(N444) );
  OAI22X1TF U594 ( .A0(N111), .A1(N1017), .B0(N502), .B1(N95), .Y(N355) );
  OAI22X1TF U595 ( .A0(N513), .A1(N512), .B0(N511), .B1(N154), .Y(N708) );
  OAI21X1TF U596 ( .A0(N507), .A1(N1008), .B0(N506), .Y(N508) );
  AOI211X1TF U597 ( .A0(SUM_AB[11]), .A1(N126), .B0(N504), .C0(N503), .Y(N506)
         );
  NAND2X2TF U598 ( .A(MODE_TYPE[1]), .B(N352), .Y(N608) );
  OAI22X1TF U599 ( .A0(N146), .A1(N89), .B0(N500), .B1(N94), .Y(N504) );
  INVX2TF U600 ( .A(N493), .Y(N507) );
  NOR2X2TF U601 ( .A(N394), .B(N1017), .Y(N493) );
  INVX2TF U602 ( .A(INTADD_0_N1), .Y(N464) );
  NOR2X1TF U603 ( .A(N151), .B(N748), .Y(INTADD_0_CI) );
  INVX2TF U604 ( .A(X_IN[0]), .Y(N748) );
  AOI31X1TF U605 ( .A0(N940), .A1(N73), .A2(N563), .B0(N349), .Y(N385) );
  OAI211X1TF U606 ( .A0(N73), .A1(N375), .B0(N359), .C0(N348), .Y(N349) );
  OAI211X1TF U607 ( .A0(N959), .A1(N347), .B0(N566), .C0(N600), .Y(N348) );
  NOR2X1TF U608 ( .A(PRE_WORK), .B(N364), .Y(N602) );
  INVX2TF U609 ( .A(N599), .Y(N566) );
  NOR2X1TF U610 ( .A(N371), .B(N943), .Y(N359) );
  INVX2TF U611 ( .A(N394), .Y(N371) );
  INVX2TF U612 ( .A(N617), .Y(N375) );
  OAI21X1TF U613 ( .A0(N759), .A1(N166), .B0(N758), .Y(N687) );
  OAI21X1TF U614 ( .A0(N757), .A1(N756), .B0(N778), .Y(N758) );
  INVX2TF U615 ( .A(N191), .Y(N778) );
  OAI211X1TF U616 ( .A0(N145), .A1(N775), .B0(N755), .C0(N754), .Y(N756) );
  AOI22X1TF U617 ( .A0(DIVISION_REMA[6]), .A1(N734), .B0(SUM_AB[7]), .B1(N136), 
        .Y(N754) );
  OAI211X1TF U618 ( .A0(N808), .A1(N996), .B0(N753), .C0(N752), .Y(N757) );
  AOI22X1TF U619 ( .A0(X_IN[1]), .A1(N805), .B0(X_IN[0]), .B1(N131), .Y(N752)
         );
  OAI21X1TF U620 ( .A0(N453), .A1(N452), .B0(N462), .Y(N996) );
  OAI22X1TF U621 ( .A0(N191), .A1(N733), .B0(N759), .B1(N164), .Y(N691) );
  AOI211X1TF U622 ( .A0(SUM_AB[3]), .A1(N137), .B0(N732), .C0(N731), .Y(N733)
         );
  OAI211X1TF U623 ( .A0(N808), .A1(N984), .B0(N755), .C0(N730), .Y(N731) );
  OAI21X1TF U624 ( .A0(N415), .A1(N414), .B0(N423), .Y(N984) );
  OAI22X1TF U625 ( .A0(N729), .A1(N802), .B0(N171), .B1(N93), .Y(N732) );
  OAI22X1TF U626 ( .A0(N191), .A1(N743), .B0(N759), .B1(N165), .Y(N689) );
  AOI211X1TF U627 ( .A0(SUM_AB[5]), .A1(N137), .B0(N742), .C0(N741), .Y(N743)
         );
  OAI211X1TF U628 ( .A0(N808), .A1(N990), .B0(N755), .C0(N740), .Y(N741) );
  AOI222X4TF U629 ( .A0(N765), .A1(N98), .B0(N763), .B1(N130), .C0(N557), .C1(
        N805), .Y(N755) );
  OAI21X1TF U630 ( .A0(N433), .A1(N432), .B0(N443), .Y(N990) );
  INVX2TF U631 ( .A(N802), .Y(N789) );
  NOR3X1TF U632 ( .A(N772), .B(N125), .C(N556), .Y(N780) );
  AOI32X1TF U633 ( .A0(N788), .A1(N814), .A2(N787), .B0(N812), .B1(N167), .Y(
        N685) );
  OAI211X1TF U634 ( .A0(N808), .A1(N1002), .B0(N784), .C0(N783), .Y(N785) );
  AOI22X1TF U635 ( .A0(DIVISION_HEAD[1]), .A1(N113), .B0(X_IN[1]), .B1(N98), 
        .Y(N783) );
  OAI21X1TF U636 ( .A0(N477), .A1(N476), .B0(N486), .Y(N1002) );
  OAI21X1TF U637 ( .A0(N782), .A1(N802), .B0(N781), .Y(N786) );
  AOI22X1TF U638 ( .A0(DIVISION_REMA[8]), .A1(N125), .B0(N798), .B1(SUM_AB[0]), 
        .Y(N781) );
  AOI22X1TF U639 ( .A0(DIVISION_HEAD[0]), .A1(N804), .B0(SUM_AB[9]), .B1(N137), 
        .Y(N788) );
  OAI21X1TF U640 ( .A0(N812), .A1(N555), .B0(N554), .Y(N706) );
  OAI21X1TF U641 ( .A0(N812), .A1(N804), .B0(DIVISION_HEAD[3]), .Y(N554) );
  AOI211X1TF U642 ( .A0(DIVISION_HEAD[2]), .A1(N125), .B0(N553), .C0(N552), 
        .Y(N555) );
  AOI22X1TF U643 ( .A0(N798), .A1(SUM_AB[3]), .B0(N1012), .B1(N795), .Y(N549)
         );
  NOR2X1TF U644 ( .A(N1017), .B(N1013), .Y(N1012) );
  AOI22X1TF U645 ( .A0(N940), .A1(SUM_AB[12]), .B0(X_IN[5]), .B1(N131), .Y(
        N550) );
  AOI22X1TF U646 ( .A0(X_IN[4]), .A1(N99), .B0(X_IN[6]), .B1(N805), .Y(N551)
         );
  OAI22X1TF U647 ( .A0(N548), .A1(N802), .B0(N547), .B1(N95), .Y(N553) );
  AOI32X1TF U648 ( .A0(N815), .A1(N814), .A2(N813), .B0(N812), .B1(N161), .Y(
        N683) );
  AOI211X1TF U649 ( .A0(DIVISION_HEAD[3]), .A1(N113), .B0(N810), .C0(N809), 
        .Y(N813) );
  OAI211X1TF U650 ( .A0(N808), .A1(N1008), .B0(N807), .C0(N806), .Y(N809) );
  AOI22X1TF U651 ( .A0(X_IN[3]), .A1(N98), .B0(X_IN[5]), .B1(N805), .Y(N806)
         );
  AND2X2TF U652 ( .A(N762), .B(N767), .Y(N764) );
  INVX2TF U653 ( .A(N386), .Y(N772) );
  AOI22X1TF U654 ( .A0(DIVISION_HEAD[1]), .A1(N125), .B0(DIVISION_HEAD[2]), 
        .B1(N804), .Y(N807) );
  INVX2TF U655 ( .A(N454), .Y(N804) );
  OAI21X1TF U656 ( .A0(N499), .A1(N498), .B0(N1013), .Y(N1008) );
  INVX2TF U657 ( .A(SUM_AB[11]), .Y(N498) );
  INVX2TF U658 ( .A(SUM_AB[9]), .Y(N476) );
  INVX2TF U659 ( .A(SUM_AB[7]), .Y(N452) );
  NOR2X1TF U660 ( .A(SUM_AB[6]), .B(N443), .Y(N453) );
  INVX2TF U661 ( .A(SUM_AB[5]), .Y(N432) );
  NOR2X1TF U662 ( .A(SUM_AB[4]), .B(N423), .Y(N433) );
  INVX2TF U663 ( .A(SUM_AB[3]), .Y(N414) );
  NOR3X1TF U664 ( .A(SUM_AB[0]), .B(SUM_AB[2]), .C(SUM_AB[1]), .Y(N415) );
  INVX2TF U665 ( .A(N795), .Y(N808) );
  NOR2X2TF U666 ( .A(N1017), .B(N649), .Y(N795) );
  INVX2TF U667 ( .A(SUM_AB[12]), .Y(N1017) );
  OAI21X1TF U668 ( .A0(N803), .A1(N802), .B0(N801), .Y(N810) );
  INVX2TF U669 ( .A(N94), .Y(N800) );
  NAND2X2TF U670 ( .A(N352), .B(N311), .Y(N802) );
  INVX2TF U671 ( .A(N812), .Y(N814) );
  INVX2TF U672 ( .A(N352), .Y(N639) );
  AOI31X1TF U673 ( .A0(N122), .A1(N384), .A2(N383), .B0(N382), .Y(N546) );
  INVX2TF U674 ( .A(N304), .Y(N763) );
  OAI211X1TF U675 ( .A0(X_IN[12]), .A1(N547), .B0(N303), .C0(N302), .Y(N304)
         );
  OAI22X1TF U676 ( .A0(Y_IN[10]), .A1(N301), .B0(N300), .B1(N299), .Y(N302) );
  OAI22X1TF U677 ( .A0(X_IN[10]), .A1(N298), .B0(X_IN[11]), .B1(N782), .Y(N299) );
  OAI21X1TF U678 ( .A0(Y_IN[9]), .A1(N297), .B0(Y_IN[8]), .Y(N298) );
  AOI211X1TF U679 ( .A0(X_IN[10]), .A1(N760), .B0(N296), .C0(N295), .Y(N300)
         );
  AOI21X1TF U680 ( .A0(Y_IN[7]), .A1(N500), .B0(N294), .Y(N295) );
  AOI211X1TF U681 ( .A0(X_IN[8]), .A1(N293), .B0(N292), .C0(N291), .Y(N294) );
  NOR2X1TF U682 ( .A(N83), .B(N500), .Y(N292) );
  AOI21X1TF U683 ( .A0(N192), .A1(N468), .B0(N290), .Y(N293) );
  AOI211X1TF U684 ( .A0(X_IN[6]), .A1(N289), .B0(N288), .C0(N287), .Y(N290) );
  NOR2X1TF U685 ( .A(N192), .B(N468), .Y(N288) );
  AOI32X1TF U686 ( .A0(N286), .A1(N285), .A2(N315), .B0(N284), .B1(N285), .Y(
        N289) );
  OAI22X1TF U687 ( .A0(X_IN[4]), .A1(N736), .B0(N100), .B1(N729), .Y(N284) );
  OAI32X1TF U688 ( .A0(N283), .A1(N84), .A2(N313), .B0(X_IN[2]), .B1(N283), 
        .Y(N286) );
  INVX2TF U689 ( .A(X_IN[7]), .Y(N468) );
  INVX2TF U690 ( .A(X_IN[9]), .Y(N500) );
  NOR2X1TF U691 ( .A(Y_IN[9]), .B(N297), .Y(N296) );
  INVX2TF U692 ( .A(X_IN[11]), .Y(N297) );
  NOR2X1TF U693 ( .A(Y_IN[12]), .B(Y_IN[11]), .Y(N303) );
  INVX2TF U694 ( .A(N768), .Y(N557) );
  OR2X2TF U695 ( .A(MODE_TYPE[0]), .B(N311), .Y(N767) );
  INVX2TF U696 ( .A(MODE_TYPE[1]), .Y(N311) );
  OAI31X1TF U697 ( .A0(N279), .A1(N278), .A2(N277), .B0(N276), .Y(N280) );
  NOR2X1TF U698 ( .A(X_IN[10]), .B(N782), .Y(N277) );
  AOI211X1TF U699 ( .A0(X_IN[10]), .A1(N782), .B0(X_IN[9]), .C0(N760), .Y(N278) );
  AOI211X1TF U700 ( .A0(X_IN[9]), .A1(N760), .B0(N275), .C0(N274), .Y(N279) );
  AOI21X1TF U701 ( .A0(Y_IN[7]), .A1(N488), .B0(N273), .Y(N274) );
  AOI211X1TF U702 ( .A0(N272), .A1(X_IN[7]), .B0(N271), .C0(N270), .Y(N273) );
  NOR2X1TF U703 ( .A(Y_IN[7]), .B(N488), .Y(N271) );
  AOI21X1TF U704 ( .A0(N192), .A1(N463), .B0(N269), .Y(N272) );
  AOI211X1TF U705 ( .A0(N268), .A1(X_IN[5]), .B0(N267), .C0(N266), .Y(N269) );
  NOR2X1TF U706 ( .A(N192), .B(N463), .Y(N267) );
  AOI211X1TF U707 ( .A0(Y_IN[3]), .A1(N442), .B0(N265), .C0(N264), .Y(N268) );
  AOI211X1TF U708 ( .A0(X_IN[4]), .A1(N729), .B0(N84), .C0(N736), .Y(N264) );
  OAI32X1TF U709 ( .A0(N263), .A1(X_IN[2]), .A2(N313), .B0(X_IN[1]), .B1(N263), 
        .Y(N265) );
  OAI211X1TF U710 ( .A0(Y_IN[3]), .A1(N442), .B0(N262), .C0(N315), .Y(N263) );
  AOI22X1TF U711 ( .A0(N84), .A1(N736), .B0(X_IN[2]), .B1(N314), .Y(N262) );
  INVX2TF U712 ( .A(X_IN[4]), .Y(N442) );
  INVX2TF U713 ( .A(X_IN[6]), .Y(N463) );
  INVX2TF U714 ( .A(X_IN[8]), .Y(N488) );
  NOR2X1TF U715 ( .A(Y_IN[9]), .B(N502), .Y(N275) );
  INVX2TF U716 ( .A(X_IN[10]), .Y(N502) );
  NOR2X1TF U717 ( .A(Y_IN[11]), .B(N301), .Y(N281) );
  INVX2TF U718 ( .A(X_IN[12]), .Y(N301) );
  INVX2TF U719 ( .A(N338), .Y(N384) );
  AOI22X1TF U720 ( .A0(N798), .A1(SUM_AB[2]), .B0(SUM_AB[11]), .B1(N137), .Y(
        N815) );
  OAI21X1TF U721 ( .A0(N170), .A1(N108), .B0(N255), .Y(OPER_A[12]) );
  INVX2TF U722 ( .A(N558), .Y(N798) );
  OAI211X1TF U723 ( .A0(N855), .A1(N854), .B0(N853), .C0(N852), .Y(N678) );
  AOI32X1TF U724 ( .A0(N936), .A1(OPER_B[4]), .A2(N851), .B0(N883), .B1(
        OPER_B[4]), .Y(N852) );
  AOI211X1TF U725 ( .A0(N857), .A1(OPER_B[5]), .B0(N850), .C0(N849), .Y(N853)
         );
  OAI31X1TF U726 ( .A0(N933), .A1(OPER_A[4]), .A2(N848), .B0(N204), .Y(N849)
         );
  AOI21X1TF U727 ( .A0(N103), .A1(C152_DATA4_4), .B0(N206), .Y(N204) );
  NOR3X1TF U728 ( .A(OPER_B[4]), .B(N851), .C(N106), .Y(N850) );
  AOI21X1TF U729 ( .A0(N930), .A1(N848), .B0(N847), .Y(N854) );
  INVX2TF U730 ( .A(N931), .Y(N847) );
  INVX2TF U731 ( .A(OPER_A[0]), .Y(N824) );
  OAI21X1TF U732 ( .A0(N152), .A1(N97), .B0(N230), .Y(FOUT[4]) );
  AOI21X1TF U733 ( .A0(N219), .A1(DIVISION_REMA[4]), .B0(N229), .Y(N230) );
  OAI22X1TF U734 ( .A0(N153), .A1(N86), .B0(N173), .B1(N80), .Y(N229) );
  AOI211X1TF U735 ( .A0(N104), .A1(C152_DATA4_5), .B0(N859), .C0(N210), .Y(
        N211) );
  OAI31X1TF U736 ( .A0(OPER_B[5]), .A1(N858), .A2(N106), .B0(N904), .Y(N859)
         );
  OAI211X1TF U737 ( .A0(SIGN_Y), .A1(N964), .B0(N220), .C0(N970), .Y(N904) );
  AOI22X1TF U738 ( .A0(N857), .A1(OPER_B[6]), .B0(N856), .B1(N861), .Y(N866)
         );
  NOR2X1TF U739 ( .A(N933), .B(OPER_A[5]), .Y(N856) );
  INVX2TF U740 ( .A(N893), .Y(N857) );
  AOI22X1TF U741 ( .A0(OPER_B[5]), .A1(N863), .B0(OPER_A[5]), .B1(N862), .Y(
        N865) );
  OAI21X1TF U742 ( .A0(N933), .A1(N861), .B0(N931), .Y(N862) );
  OAI21X1TF U743 ( .A0(N106), .A1(N860), .B0(N934), .Y(N863) );
  OAI21X1TF U744 ( .A0(N142), .A1(N96), .B0(N224), .Y(FOUT[1]) );
  AOI21X1TF U745 ( .A0(N219), .A1(DIVISION_REMA[1]), .B0(N223), .Y(N224) );
  OAI22X1TF U746 ( .A0(N143), .A1(N85), .B0(N164), .B1(N79), .Y(N223) );
  OAI211X1TF U747 ( .A0(N893), .A1(N159), .B0(N892), .C0(N891), .Y(N675) );
  AOI211X1TF U748 ( .A0(OPER_A[7]), .A1(N889), .B0(N888), .C0(N887), .Y(N892)
         );
  INVX2TF U749 ( .A(N207), .Y(N887) );
  AOI211X1TF U750 ( .A0(N103), .A1(C152_DATA4_7), .B0(N206), .C0(N205), .Y(
        N207) );
  NOR3X1TF U751 ( .A(N105), .B(OPER_B[7]), .C(N886), .Y(N205) );
  OR2X2TF U752 ( .A(N929), .B(N885), .Y(N206) );
  NOR2X1TF U753 ( .A(N966), .B(N829), .Y(N869) );
  INVX2TF U754 ( .A(N884), .Y(N888) );
  AOI32X1TF U755 ( .A0(OPER_B[7]), .A1(N936), .A2(N886), .B0(N883), .B1(
        OPER_B[7]), .Y(N884) );
  INVX2TF U756 ( .A(N934), .Y(N883) );
  OAI21X1TF U757 ( .A0(N933), .A1(N890), .B0(N931), .Y(N889) );
  NOR3X1TF U758 ( .A(N73), .B(N177), .C(N964), .Y(N963) );
  OAI22X1TF U759 ( .A0(N189), .A1(N200), .B0(N201), .B1(OFFSET[2]), .Y(C2_Z_4)
         );
  INVX2TF U760 ( .A(Y_IN[4]), .Y(N200) );
  OAI22X1TF U761 ( .A0(N189), .A1(N199), .B0(N201), .B1(OFFSET[3]), .Y(C2_Z_5)
         );
  OAI22X1TF U762 ( .A0(N189), .A1(N198), .B0(N201), .B1(OFFSET[4]), .Y(C2_Z_6)
         );
  OAI22X1TF U763 ( .A0(N189), .A1(N193), .B0(N201), .B1(OFFSET[5]), .Y(C2_Z_7)
         );
  OAI22X1TF U764 ( .A0(N189), .A1(N760), .B0(N201), .B1(OFFSET[6]), .Y(C2_Z_8)
         );
  OAI22X1TF U765 ( .A0(N189), .A1(N782), .B0(N201), .B1(OFFSET[7]), .Y(C2_Z_9)
         );
  OAI22X1TF U766 ( .A0(N189), .A1(N547), .B0(N132), .B1(OFFSET[8]), .Y(C2_Z_10) );
  OAI22X1TF U767 ( .A0(N189), .A1(N803), .B0(N132), .B1(OFFSET[9]), .Y(C2_Z_11) );
  INVX2TF U768 ( .A(Y_IN[11]), .Y(N803) );
  NOR2X1TF U769 ( .A(OPER_B[9]), .B(N907), .Y(N922) );
  NOR2X1TF U770 ( .A(N868), .B(OPER_B[6]), .Y(N886) );
  INVX2TF U771 ( .A(N872), .Y(N868) );
  NOR2X1TF U772 ( .A(OPER_B[5]), .B(N860), .Y(N872) );
  NOR2X1TF U773 ( .A(OPER_B[3]), .B(N840), .Y(N851) );
  AOI211X1TF U774 ( .A0(N56), .A1(N964), .B0(SIGN_Y), .C0(N909), .Y(N929) );
  NOR2X1TF U775 ( .A(OPER_A[9]), .B(N908), .Y(N916) );
  NOR2X1TF U776 ( .A(OPER_A[7]), .B(N890), .Y(N897) );
  NOR2X1TF U777 ( .A(OPER_A[5]), .B(N861), .Y(N875) );
  NOR2X1TF U778 ( .A(OPER_A[3]), .B(N839), .Y(N848) );
  OAI21X1TF U779 ( .A0(N152), .A1(N108), .B0(N246), .Y(OPER_A[4]) );
  OAI21X1TF U780 ( .A0(N144), .A1(N108), .B0(N247), .Y(OPER_A[5]) );
  OAI21X1TF U781 ( .A0(N153), .A1(N108), .B0(N248), .Y(OPER_A[6]) );
  OAI21X1TF U782 ( .A0(N141), .A1(N108), .B0(N249), .Y(OPER_A[7]) );
  OAI21X1TF U783 ( .A0(N175), .A1(N108), .B0(N250), .Y(OPER_A[8]) );
  OAI21X1TF U784 ( .A0(N108), .A1(N528), .B0(N251), .Y(OPER_A[9]) );
  OAI21X1TF U785 ( .A0(N108), .A1(N146), .B0(N252), .Y(OPER_A[10]) );
  OAI21X1TF U786 ( .A0(N108), .A1(N154), .B0(N253), .Y(OPER_A[11]) );
  OAI211X1TF U787 ( .A0(N176), .A1(N937), .B0(N846), .C0(N845), .Y(N679) );
  AOI211X1TF U788 ( .A0(OPER_A[3]), .A1(N844), .B0(N843), .C0(N842), .Y(N845)
         );
  OAI31X1TF U789 ( .A0(N933), .A1(OPER_A[3]), .A2(N841), .B0(N203), .Y(N842)
         );
  AOI21X1TF U790 ( .A0(C152_DATA4_3), .A1(N103), .B0(N905), .Y(N203) );
  OAI22X1TF U791 ( .A0(N969), .A1(N729), .B0(N201), .B1(OFFSET[1]), .Y(C2_Z_3)
         );
  INVX2TF U792 ( .A(DP_OP_333_124_4748_N57), .Y(N201) );
  INVX2TF U793 ( .A(Y_IN[3]), .Y(N729) );
  OAI32X1TF U794 ( .A0(N182), .A1(N105), .A2(N840), .B0(N934), .B1(N182), .Y(
        N843) );
  INVX2TF U795 ( .A(N867), .Y(N920) );
  AOI32X1TF U796 ( .A0(N605), .A1(N346), .A2(N822), .B0(N945), .B1(N345), .Y(
        N867) );
  INVX2TF U797 ( .A(N939), .Y(N945) );
  OAI21X1TF U798 ( .A0(N933), .A1(N839), .B0(N931), .Y(N844) );
  INVX2TF U799 ( .A(N830), .Y(N911) );
  AOI21X1TF U800 ( .A0(N564), .A1(N345), .B0(N563), .Y(N830) );
  INVX2TF U801 ( .A(N841), .Y(N839) );
  NOR3X1TF U802 ( .A(OPER_A[2]), .B(OPER_A[1]), .C(OPER_A[0]), .Y(N841) );
  OAI21X1TF U803 ( .A0(N150), .A1(N107), .B0(N244), .Y(OPER_A[2]) );
  INVX2TF U804 ( .A(N930), .Y(N933) );
  NOR2X2TF U805 ( .A(N923), .B(N915), .Y(N930) );
  INVX2TF U806 ( .A(N903), .Y(N923) );
  OAI21X1TF U807 ( .A0(N143), .A1(N107), .B0(N245), .Y(OPER_A[3]) );
  AOI31X1TF U808 ( .A0(N936), .A1(N182), .A2(N840), .B0(N881), .Y(N846) );
  OAI21X1TF U809 ( .A0(N974), .A1(N909), .B0(N836), .Y(N881) );
  INVX2TF U810 ( .A(N909), .Y(N220) );
  INVX2TF U811 ( .A(N344), .Y(N958) );
  INVX2TF U812 ( .A(N565), .Y(N948) );
  NOR2X1TF U813 ( .A(OPER_B[1]), .B(OPER_B[0]), .Y(N832) );
  INVX2TF U814 ( .A(N345), .Y(N346) );
  INVX2TF U815 ( .A(N605), .Y(N821) );
  NOR2X2TF U816 ( .A(N603), .B(N631), .Y(N822) );
  AOI221X1TF U817 ( .A0(N128), .A1(N157), .B0(N180), .B1(N91), .C0(N817), .Y(
        N818) );
  AOI22X1TF U818 ( .A0(\INDEX[2] ), .A1(N90), .B0(N124), .B1(\RSHT_BITS[3] ), 
        .Y(N816) );
  AOI32X1TF U819 ( .A0(N939), .A1(N952), .A2(N368), .B0(N954), .B1(N952), .Y(
        N342) );
  OR2X2TF U820 ( .A(N631), .B(N148), .Y(N368) );
  INVX2TF U821 ( .A(N603), .Y(N642) );
  OAI21X1TF U822 ( .A0(N344), .A1(N938), .B0(N340), .Y(N607) );
  OAI21X1TF U823 ( .A0(N570), .A1(N564), .B0(N341), .Y(N340) );
  NOR2X2TF U824 ( .A(\RSHT_BITS[3] ), .B(N591), .Y(N605) );
  NOR3X1TF U825 ( .A(N121), .B(N122), .C(N953), .Y(N820) );
  INVX2TF U826 ( .A(N959), .Y(N966) );
  NOR2X1TF U827 ( .A(SIGN_Y), .B(N109), .Y(N906) );
  INVX2TF U828 ( .A(N308), .Y(N627) );
  OAI22X1TF U829 ( .A0(Y_IN[12]), .A1(N175), .B0(N336), .B1(N335), .Y(N337) );
  OAI31X1TF U830 ( .A0(N334), .A1(DIVISION_HEAD[10]), .A2(N547), .B0(N333), 
        .Y(N335) );
  AOI22X1TF U831 ( .A0(Y_IN[11]), .A1(N141), .B0(N332), .B1(N331), .Y(N333) );
  OAI22X1TF U832 ( .A0(DIVISION_HEAD[8]), .A1(N760), .B0(DIVISION_HEAD[9]), 
        .B1(N782), .Y(N331) );
  INVX2TF U833 ( .A(N330), .Y(N332) );
  NOR2X1TF U834 ( .A(Y_IN[11]), .B(N141), .Y(N334) );
  AOI211X1TF U835 ( .A0(DIVISION_HEAD[8]), .A1(N760), .B0(N329), .C0(N330), 
        .Y(N336) );
  OAI21X1TF U836 ( .A0(Y_IN[11]), .A1(N141), .B0(N328), .Y(N330) );
  AOI22X1TF U837 ( .A0(DIVISION_HEAD[10]), .A1(N547), .B0(DIVISION_HEAD[9]), 
        .B1(N782), .Y(N328) );
  INVX2TF U838 ( .A(Y_IN[9]), .Y(N782) );
  INVX2TF U839 ( .A(Y_IN[10]), .Y(N547) );
  AOI21X1TF U840 ( .A0(N83), .A1(N143), .B0(N327), .Y(N329) );
  AOI211X1TF U841 ( .A0(N326), .A1(DIVISION_HEAD[6]), .B0(N325), .C0(N324), 
        .Y(N327) );
  NOR2X1TF U842 ( .A(N83), .B(N143), .Y(N325) );
  AOI21X1TF U843 ( .A0(N192), .A1(N142), .B0(N323), .Y(N326) );
  AOI211X1TF U844 ( .A0(N322), .A1(DIVISION_HEAD[4]), .B0(N321), .C0(N320), 
        .Y(N323) );
  NOR2X1TF U845 ( .A(Y_IN[5]), .B(N142), .Y(N321) );
  AOI21X1TF U846 ( .A0(Y_IN[3]), .A1(N147), .B0(N319), .Y(N322) );
  OAI32X1TF U847 ( .A0(N318), .A1(DIVISION_HEAD[2]), .A2(N736), .B0(N317), 
        .B1(N318), .Y(N319) );
  OAI211X1TF U848 ( .A0(Y_IN[2]), .A1(N161), .B0(N316), .C0(N315), .Y(N317) );
  INVX2TF U849 ( .A(Y_IN[0]), .Y(N655) );
  INVX2TF U850 ( .A(Y_IN[1]), .Y(N313) );
  INVX2TF U851 ( .A(Y_IN[2]), .Y(N736) );
  NOR2X1TF U852 ( .A(Y_IN[3]), .B(N147), .Y(N318) );
  INVX2TF U853 ( .A(Y_IN[8]), .Y(N760) );
  INVX2TF U854 ( .A(Y_IN[12]), .Y(N548) );
  OAI21X1TF U855 ( .A0(N175), .A1(N97), .B0(N238), .Y(FOUT[8]) );
  AOI21X1TF U856 ( .A0(N219), .A1(DIVISION_REMA[8]), .B0(N237), .Y(N238) );
  OAI22X1TF U857 ( .A0(N172), .A1(N80), .B0(N146), .B1(N85), .Y(N237) );
  OAI21X1TF U858 ( .A0(N144), .A1(N96), .B0(N232), .Y(FOUT[5]) );
  AOI21X1TF U859 ( .A0(N219), .A1(DIVISION_REMA[5]), .B0(N231), .Y(N232) );
  OAI22X1TF U860 ( .A0(N141), .A1(N85), .B0(N166), .B1(N79), .Y(N231) );
  OAI21X1TF U861 ( .A0(N141), .A1(N97), .B0(N236), .Y(FOUT[7]) );
  AOI21X1TF U862 ( .A0(N219), .A1(DIVISION_REMA[7]), .B0(N235), .Y(N236) );
  OAI22X1TF U863 ( .A0(N167), .A1(N80), .B0(N528), .B1(N86), .Y(N235) );
  OAI21X1TF U864 ( .A0(N143), .A1(N96), .B0(N228), .Y(FOUT[3]) );
  AOI21X1TF U865 ( .A0(N219), .A1(DIVISION_REMA[3]), .B0(N227), .Y(N228) );
  OAI22X1TF U866 ( .A0(N144), .A1(N85), .B0(N165), .B1(N79), .Y(N227) );
  OAI21X1TF U867 ( .A0(N153), .A1(N97), .B0(N234), .Y(FOUT[6]) );
  AOI21X1TF U868 ( .A0(N219), .A1(DIVISION_REMA[6]), .B0(N233), .Y(N234) );
  OAI22X1TF U869 ( .A0(N175), .A1(N86), .B0(N145), .B1(N79), .Y(N233) );
  OAI21X1TF U870 ( .A0(N150), .A1(N96), .B0(N226), .Y(FOUT[2]) );
  AOI21X1TF U871 ( .A0(N219), .A1(DIVISION_REMA[2]), .B0(N225), .Y(N226) );
  OAI22X1TF U872 ( .A0(N152), .A1(N85), .B0(N168), .B1(N79), .Y(N225) );
  NOR2X1TF U873 ( .A(N338), .B(N369), .Y(ALU_IS_DONE) );
  OAI211X1TF U874 ( .A0(N150), .A1(N86), .B0(N222), .C0(N221), .Y(FOUT[0]) );
  AOI22X1TF U875 ( .A0(N118), .A1(\INTADD_0_SUM[5] ), .B0(N798), .B1(
        SUM_AB[10]), .Y(N448) );
  AOI21X1TF U876 ( .A0(N118), .A1(N472), .B0(N471), .Y(N473) );
  AOI22X1TF U877 ( .A0(N117), .A1(N465), .B0(SUM_AB[8]), .B1(N126), .Y(N467)
         );
  AOI22X1TF U878 ( .A0(N118), .A1(\INTADD_0_SUM[3] ), .B0(SUM_AB[4]), .B1(N127), .Y(N431) );
  AOI31X1TF U879 ( .A0(X_IN[0]), .A1(N118), .A2(N151), .B0(N390), .Y(N391) );
  AOI22X1TF U880 ( .A0(N118), .A1(\INTADD_0_SUM[1] ), .B0(SUM_AB[2]), .B1(N127), .Y(N412) );
  AOI22X1TF U881 ( .A0(N118), .A1(\INTADD_0_SUM[0] ), .B0(SUM_AB[1]), .B1(N127), .Y(N402) );
  AOI22X1TF U882 ( .A0(N118), .A1(\INTADD_0_SUM[6] ), .B0(SUM_AB[7]), .B1(N127), .Y(N461) );
  AOI31X1TF U883 ( .A0(N117), .A1(N146), .A2(N494), .B0(N489), .Y(N490) );
  AOI22X1TF U884 ( .A0(N117), .A1(\INTADD_0_SUM[4] ), .B0(SUM_AB[5]), .B1(N126), .Y(N438) );
  AOI22X1TF U885 ( .A0(N118), .A1(\INTADD_0_SUM[2] ), .B0(SUM_AB[3]), .B1(N127), .Y(N422) );
  AOI21X1TF U886 ( .A0(N118), .A1(N356), .B0(N513), .Y(N357) );
  AOI31X1TF U887 ( .A0(N118), .A1(N154), .A2(N510), .B0(N508), .Y(N512) );
  NOR2X1TF U888 ( .A(ALU_TYPE[2]), .B(ALU_TYPE[0]), .Y(N196) );
  NAND3X1TF U889 ( .A(N904), .B(N214), .C(N213), .Y(N674) );
  NAND4BX1TF U890 ( .AN(N837), .B(N209), .C(N838), .D(N208), .Y(N680) );
  AOI2BB2X1TF U891 ( .B0(N104), .B1(C152_DATA4_2), .A0N(N155), .A1N(N928), .Y(
        N208) );
  OAI2BB1X1TF U892 ( .A0N(N104), .A1N(C152_DATA4_10), .B0(N215), .Y(N672) );
  NAND3X1TF U893 ( .A(N865), .B(N866), .C(N211), .Y(N677) );
  OAI2BB2XLTF U894 ( .B0(OFFSET[0]), .B1(N201), .A0N(Y_IN[2]), .A1N(N120), .Y(
        C2_Z_2) );
  AOI2BB2X1TF U895 ( .B0(N219), .B1(DIVISION_REMA[0]), .A0N(N171), .A1N(N80), 
        .Y(N222) );
  OAI222X1TF U896 ( .A0(N96), .A1(N528), .B0(N80), .B1(N161), .C0(N154), .C1(
        N86), .Y(FOUT[9]) );
  NAND2X1TF U897 ( .A(N148), .B(N163), .Y(N369) );
  NAND3X1TF U898 ( .A(STEP[2]), .B(STEP[3]), .C(N642), .Y(N939) );
  NAND3X1TF U899 ( .A(N545), .B(N386), .C(N634), .Y(N647) );
  NOR4XLTF U900 ( .A(N761), .B(N617), .C(N800), .D(N647), .Y(N261) );
  AOI222XLTF U901 ( .A0(STEP[2]), .A1(N149), .B0(N121), .B1(N163), .C0(N140), 
        .C1(N122), .Y(N259) );
  NAND3X1TF U902 ( .A(N261), .B(N360), .C(N633), .Y(N619) );
  AOI2BB1X1TF U903 ( .A0N(X_IN[5]), .A1N(N268), .B0(Y_IN[4]), .Y(N266) );
  AOI2BB1X1TF U904 ( .A0N(X_IN[7]), .A1N(N272), .B0(Y_IN[6]), .Y(N270) );
  NAND2X1TF U905 ( .A(MODE_TYPE[0]), .B(N311), .Y(N762) );
  AO22X1TF U906 ( .A0(X_IN[4]), .A1(N736), .B0(N84), .B1(N314), .Y(N283) );
  NAND2X1TF U907 ( .A(N100), .B(N729), .Y(N285) );
  AOI2BB1X1TF U908 ( .A0N(N289), .A1N(X_IN[6]), .B0(Y_IN[4]), .Y(N287) );
  AOI2BB1X1TF U909 ( .A0N(N293), .A1N(X_IN[8]), .B0(Y_IN[6]), .Y(N291) );
  NAND2X1TF U910 ( .A(N156), .B(N180), .Y(N616) );
  NAND4BX1TF U911 ( .AN(N382), .B(N312), .C(N802), .D(N360), .Y(N725) );
  NAND2X1TF U912 ( .A(N832), .B(N155), .Y(N840) );
  NAND2X1TF U913 ( .A(N851), .B(N176), .Y(N860) );
  NOR2BX1TF U914 ( .AN(N886), .B(OPER_B[7]), .Y(N894) );
  NAND2X1TF U915 ( .A(N894), .B(N159), .Y(N907) );
  NAND2X1TF U916 ( .A(N922), .B(N160), .Y(N935) );
  NAND2X1TF U917 ( .A(N906), .B(N74), .Y(N957) );
  NAND2X1TF U918 ( .A(N565), .B(N957), .Y(N938) );
  NAND2X1TF U919 ( .A(N966), .B(N377), .Y(N573) );
  NAND3X1TF U920 ( .A(N92), .B(N91), .C(N90), .Y(N591) );
  NOR2BX1TF U921 ( .AN(N573), .B(N605), .Y(N570) );
  NAND2X1TF U922 ( .A(PRE_WORK), .B(N350), .Y(N952) );
  NAND2X1TF U923 ( .A(N605), .B(N822), .Y(N343) );
  NAND2X1TF U924 ( .A(N218), .B(N958), .Y(N362) );
  NAND3X1TF U925 ( .A(SIGN_Y), .B(N74), .C(N905), .Y(N823) );
  NAND2X1TF U926 ( .A(N855), .B(N848), .Y(N861) );
  NAND2X1TF U927 ( .A(N874), .B(N875), .Y(N890) );
  NAND2X1TF U928 ( .A(N896), .B(N897), .Y(N908) );
  NAND2X1TF U929 ( .A(N914), .B(N916), .Y(N932) );
  NAND3X1TF U930 ( .A(N605), .B(N602), .C(N162), .Y(N600) );
  NAND2X1TF U931 ( .A(N415), .B(N414), .Y(N423) );
  NAND2X1TF U932 ( .A(N433), .B(N432), .Y(N443) );
  NAND2X1TF U933 ( .A(N453), .B(N452), .Y(N462) );
  NAND2X1TF U934 ( .A(N499), .B(N498), .Y(N1013) );
  AOI222XLTF U935 ( .A0(XTEMP[11]), .A1(X_IN[11]), .B0(XTEMP[11]), .B1(N497), 
        .C0(X_IN[11]), .C1(N497), .Y(N351) );
  XOR2X1TF U936 ( .A(X_IN[12]), .B(N351), .Y(N356) );
  NAND3X1TF U937 ( .A(N566), .B(POST_WORK), .C(N602), .Y(N372) );
  NAND3BX1TF U938 ( .AN(N362), .B(N948), .C(N966), .Y(N598) );
  NAND3X1TF U939 ( .A(N609), .B(N363), .C(N598), .Y(N942) );
  NAND2X1TF U940 ( .A(N111), .B(N394), .Y(N381) );
  NAND3X1TF U941 ( .A(N384), .B(N122), .C(DP_OP_333_124_4748_N57), .Y(N638) );
  NOR2BX1TF U942 ( .AN(N634), .B(N943), .Y(N542) );
  NAND3X1TF U943 ( .A(N542), .B(N376), .C(N375), .Y(N380) );
  NAND4X1TF U944 ( .A(N427), .B(N426), .C(N425), .D(N424), .Y(N428) );
  NAND4X1TF U945 ( .A(N438), .B(N437), .C(N436), .D(N435), .Y(N439) );
  NAND4X1TF U946 ( .A(N448), .B(N447), .C(N446), .D(N445), .Y(N449) );
  OAI2BB1X1TF U947 ( .A0N(DIVISION_HEAD[10]), .A1N(N471), .B0(N451), .Y(N713)
         );
  AOI2BB2X1TF U948 ( .B0(X_IN[9]), .B1(N478), .A0N(N478), .A1N(X_IN[9]), .Y(
        N483) );
  NAND3X1TF U949 ( .A(N117), .B(N528), .C(N483), .Y(N479) );
  AOI2BB1X1TF U950 ( .A0N(N509), .A1N(N483), .B0(N513), .Y(N484) );
  AOI2BB2X1TF U951 ( .B0(N487), .B1(N502), .A0N(N502), .A1N(N487), .Y(N494) );
  AOI2BB1X1TF U952 ( .A0N(N509), .A1N(N494), .B0(N513), .Y(N495) );
  AOI2BB2X1TF U953 ( .B0(N78), .B1(N497), .A0N(N497), .A1N(N78), .Y(N510) );
  OAI2BB2XLTF U954 ( .B0(N502), .B1(N608), .A0N(XTEMP[12]), .A1N(N87), .Y(N503) );
  AOI2BB1X1TF U955 ( .A0N(N509), .A1N(N510), .B0(N513), .Y(N511) );
  AOI2BB1X1TF U956 ( .A0N(DIVISION_REMA[2]), .A1N(N517), .B0(DIVISION_HEAD[6]), 
        .Y(N515) );
  OA21XLTF U957 ( .A0(N152), .A1(DIVISION_REMA[4]), .B0(N519), .Y(N521) );
  OA21XLTF U958 ( .A0(N153), .A1(DIVISION_REMA[6]), .B0(N523), .Y(N525) );
  OA21XLTF U959 ( .A0(XTEMP[12]), .A1(N535), .B0(N147), .Y(N534) );
  NAND4X1TF U960 ( .A(N545), .B(N544), .C(N638), .D(N543), .Y(N556) );
  NAND3X1TF U961 ( .A(N551), .B(N550), .C(N549), .Y(N552) );
  NAND3X1TF U962 ( .A(N755), .B(N559), .C(N558), .Y(N560) );
  NAND3X1TF U963 ( .A(N566), .B(N602), .C(N821), .Y(N572) );
  NAND4X1TF U964 ( .A(N568), .B(N567), .C(N639), .D(N572), .Y(N569) );
  NAND2X1TF U965 ( .A(N179), .B(N157), .Y(N590) );
  NOR4XLTF U966 ( .A(\RSHT_BITS[3] ), .B(N90), .C(N614), .D(N590), .Y(N571) );
  NAND2X1TF U967 ( .A(N579), .B(N589), .Y(N586) );
  NAND2X1TF U968 ( .A(N92), .B(N91), .Y(N588) );
  AOI2BB2X1TF U969 ( .B0(N596), .B1(N157), .A0N(N590), .A1N(N592), .Y(N584) );
  NAND4X1TF U970 ( .A(N93), .B(N634), .C(N633), .D(N632), .Y(N635) );
  NAND4X1TF U971 ( .A(N640), .B(N639), .C(N638), .D(N643), .Y(N697) );
  NAND3X1TF U972 ( .A(N755), .B(N651), .C(N650), .Y(N652) );
  AO22X1TF U973 ( .A0(DIVISION_REMA[4]), .A1(N734), .B0(N192), .B1(N789), .Y(
        N742) );
  AOI2BB1X1TF U974 ( .A0N(X_IN[1]), .A1N(N763), .B0(N762), .Y(N766) );
  NAND4X1TF U975 ( .A(N793), .B(N792), .C(N791), .D(N790), .Y(N794) );
  OAI221XLTF U976 ( .A0(\INDEX[2] ), .A1(N90), .B0(N124), .B1(\RSHT_BITS[3] ), 
        .C0(N816), .Y(N817) );
  OAI221XLTF U977 ( .A0(N129), .A1(N179), .B0(N156), .B1(N92), .C0(N818), .Y(
        N829) );
  NAND2X1TF U978 ( .A(N903), .B(N869), .Y(N864) );
  NAND2BX1TF U979 ( .AN(N819), .B(N864), .Y(N885) );
  NAND2X1TF U980 ( .A(N828), .B(N966), .Y(N870) );
  NAND3X1TF U981 ( .A(SIGN_Y), .B(N74), .C(N220), .Y(N836) );
  OAI2BB1X1TF U982 ( .A0N(N959), .A1N(N829), .B0(N828), .Y(N919) );
  NAND3X1TF U983 ( .A(N74), .B(N177), .C(N56), .Y(N974) );
  NAND4X1TF U984 ( .A(N220), .B(N177), .C(N56), .D(N964), .Y(N838) );
  NAND2X1TF U985 ( .A(N903), .B(N919), .Y(N937) );
  NAND3BX1TF U986 ( .AN(OPER_A[7]), .B(N930), .C(N890), .Y(N891) );
  NAND2X1TF U987 ( .A(N940), .B(N945), .Y(N946) );
  NAND2X1TF U988 ( .A(N978), .B(N977), .Y(N668) );
  NAND2X1TF U989 ( .A(N981), .B(N980), .Y(N667) );
  NAND2X1TF U990 ( .A(SUM_AB[3]), .B(N82), .Y(N982) );
  NAND2X1TF U991 ( .A(N987), .B(N986), .Y(N665) );
  NAND2X1TF U992 ( .A(SUM_AB[5]), .B(N82), .Y(N988) );
  NAND2X1TF U993 ( .A(N993), .B(N992), .Y(N663) );
  NAND2X1TF U994 ( .A(SUM_AB[7]), .B(N82), .Y(N994) );
  NAND2X1TF U995 ( .A(N999), .B(N998), .Y(N661) );
  NAND2X1TF U996 ( .A(SUM_AB[9]), .B(N82), .Y(N1000) );
  NAND2X1TF U997 ( .A(N1005), .B(N1004), .Y(N659) );
  NAND2X1TF U998 ( .A(SUM_AB[11]), .B(N82), .Y(N1006) );
endmodule


module SERIAL_CPU_8BIT_VG ( CLK, ENABLE, RST_N, START, I_DATAIN, D_DATAIN, 
        IS_I_ADDR, NXT, I_ADDR, D_ADDR, D_WE, D_DATAOUT, IO_STATUS, IO_CONTROL, 
        IO_DATAINA, IO_DATAINB, IO_DATAOUTA, IO_DATAOUTB, IO_OFFSET );
  input [7:0] I_DATAIN;
  input [7:0] D_DATAIN;
  output [1:0] NXT;
  output [8:0] I_ADDR;
  output [8:0] D_ADDR;
  output [7:0] D_DATAOUT;
  input [15:0] IO_STATUS;
  output [15:0] IO_CONTROL;
  input [15:0] IO_DATAINA;
  input [15:0] IO_DATAINB;
  output [15:0] IO_DATAOUTA;
  output [15:0] IO_DATAOUTB;
  output [15:0] IO_OFFSET;
  input CLK, ENABLE, RST_N, START;
  output IS_I_ADDR, D_WE;
  wire   \OPER1_R1[2] , N110, N166, N167, N168, CF_BUF, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N504, N505, N506, N507, N508, N509, N510, N511, N512,
         N513, N514, N515, N516, N517, N518, N519, N588, N589, ZF, CF, N616,
         N400, N401, N402, N403, N404, N405, N406, N408, N409, N411, N412,
         N413, N414, N415, N416, N418, N420, N421, N423, N424, N433, N434,
         N435, N436, N437, N438, N439, N440, N441, N442, N443, N444, N445,
         N447, N448, N449, N451, N452, N453, N455, N456, N457, N459, N460,
         N461, N462, N464, N465, N466, N468, N469, N4700, N4720, N4730, N4740,
         N4750, N4770, N4780, N4790, N4800, N4820, N4830, N4840, N4860, N487,
         N488, N489, N491, N492, N493, N495, N496, N497, N498, N500, N501,
         N502, N503, N5050, N5060, N5070, N5080, N5100, N5110, N5130, N5140,
         N5180, N520, N521, N522, N523, N524, N525, N526, N527, N528, N529,
         N530, N531, N532, N533, N534, N535, N554, N569, N571, N572, N595,
         N596, N597, N598, N599, N600, N601, N602, N603, N604, N605, N606,
         N607, N608, N609, N610, N613, N614, N615, N6160, N617, N618, N619,
         N620, N621, N622, N623, N624, N625, N626, N627, N628, N629, N630,
         N631, N632, N633, N634, N635, N636, N637, N638, N639, N640, N641,
         N642, N643, N644, N645, N646, N647, N648, N649, N650, N651, N652,
         N653, N654, N655, N656, N657, N658, N659, N660, N661, N662, N663,
         N664, N665, N666, N667, N668, N669, N670, N671, N672, N673, N674,
         N675, N676, N677, N678, N679, N680, N681, N682, N683, N684, N685,
         N686, N687, N688, N689, N690, N691, N692, N804, N808, N809, N810,
         N811, N812, N859, N860, N922, N923, N924, N925, N926, N927, N928,
         N929, N930, N931, N932, N933, N934, N935, N936, N937, N938, N939,
         N940, N941, N942, N943, N944, N945, N946, N947, N948, N949, N950,
         N951, N952, N953, N954, N955, N956, N957, N958, N959, N960, N961,
         N962, N963, N964, N965, N966, N967, N968, N969, N970, N971, N972,
         N973, N974, N975, N976, N977, N978, N979, N980, N981, N982, N983,
         N984, N985, N986, N987, N988, N989, N990, N991, N992, N993, N994,
         N995, N996, N997, N998, N999, N1000, N1001, N1002, SUB_X_285_4_N16,
         SUB_X_285_4_N15, SUB_X_285_4_N14, SUB_X_285_4_N13, SUB_X_285_4_N12,
         SUB_X_285_4_N11, SUB_X_285_4_N10, SUB_X_285_4_N9, SUB_X_285_4_N8,
         SUB_X_285_4_N7, SUB_X_285_4_N6, SUB_X_285_4_N5, SUB_X_285_4_N4,
         SUB_X_285_4_N3, SUB_X_285_4_N2, SUB_X_285_4_N1, ADD_X_285_3_N16,
         ADD_X_285_3_N15, ADD_X_285_3_N14, ADD_X_285_3_N13, ADD_X_285_3_N12,
         ADD_X_285_3_N11, ADD_X_285_3_N10, ADD_X_285_3_N9, ADD_X_285_3_N8,
         ADD_X_285_3_N7, ADD_X_285_3_N6, ADD_X_285_3_N5, ADD_X_285_3_N4,
         ADD_X_285_3_N3, ADD_X_285_3_N2, N1, N2, N3, N4, N5, N6, N7, N8, N9,
         N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23,
         N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, N53, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N1660, N1670, N1680, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, N192, N193, N200, N201, N202, N203, N204,
         N205, N206, N207, N208, N209, N210, N211, N212, N213, N214, N215,
         N216, N217, N218, N219, N220, N221, N222, N223, N224, N225, N226,
         N227, N228, N229, N230, N231, N232, N233, N234, N235, N236, N237,
         N238, N239, N240, N241, N242, N243, N244, N245, N246, N247, N248,
         N249, N250, N251, N252, N253, N254, N255, N256, N257, N258, N259,
         N260, N261, N262, N263, N264, N265, N266, N267, N268, N269, N270,
         N271, N272, N273, N274, N275, N276, N277, N278, N279, N280, N281,
         N282, N283, N284, N285, N286, N287, N288, N289, N290, N291, N292,
         N293, N294, N295, N296, N297, N298, N299, N300, N301, N302, N303,
         N304, N305, N306, N307, N308, N309, N310, N311, N312, N313, N314,
         N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325,
         N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336,
         N337, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347,
         N348, N349, N350, N351, N352, N353, N354, N355, N356, N357, N358,
         N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, N369,
         N370, N371, N372, N373, N374, N375, N376, N377, N378, N379, N380,
         N381, N382, N383, N384, N385, N386, N387, N388, N389, N390, N391,
         N392, N393, N394, N395, N396, N397, N398, N399, N407, N410, N417,
         N419, N422, N425, N426, N427, N428, N429, N430, N431, N432, N446,
         N450, N454, N458, N463, N467, N4710, N4760, N4810, N4850, N490, N494,
         N499, N5040, N5090, N5120, N5150, N5160, N5170, N5190, N536, N537,
         N538, N539, N540, N541, N542, N543, N544, N545, N546, N547, N548,
         N549, N550, N551, N552, N553, N555, N556, N557, N558, N559, N560,
         N561, N562, N563, N564, N565, N566, N567, N568, N570, N573, N574,
         N575, N576, N577, N578, N579, N580, N581, N582, N583, N584, N585,
         N586, N587, N5880, N5890, N590, N591, N592, N593, N594, N611, N612,
         N693, N694, N695, N696, N697, N698, N699, N700, N701, N702, N703,
         N704, N705, N706, N707, N708, N709, N710, N711, N712, N713, N714,
         N715, N716, N717, N718, N719, N720, N721, N722, N723, N724, N725,
         N726, N727, N728, N729, N730, N731, N732, N733, N734, N735, N736,
         N737, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747,
         N748, N749, N750, N751, N752, N753, N754, N755, N756, N757, N758,
         N759, N760, N761, N762, N763, N764, N765, N766, N767, N768, N769,
         N770, N771, N772, N773, N774, N775, N776, N777, N778, N779, N780,
         N781, N782, N783, N784, N785, N786, N787, N788, N789, N790, N791,
         N792, N793, N794, N795, N796, N797, N798, N799, N800, N801, N802,
         N803, N805, N806, N807, N813, N814, N815, N816, N817, N818, N819,
         N820, N821, N822, N823, N824, N825, N826, N827, N828, N829, N830,
         N831, N832, N833, N834, N835, N836, N837, N838, N839, N840, N841,
         N842, N843, N844, N845, N846, N847, N848, N849, N850, N851, N852,
         N853, N854, N855, N856, N857, N858, N861, N862, N863, N864, N865,
         N866, N867, N868, N869, N870, N871, N872, N873, N874, N875, N876,
         N877, N878, N879, N880, N881, N882, N883, N884, N885, N886, N887,
         N888, N889, N890, N891, N892, N893, N894, N895, N896, N897, N898,
         N899, N900, N901, N902, N903, N904, N905, N906, N907, N908, N909,
         N910, N911, N912, N913, N914, N915, N916, N917, N918, N919, N920,
         N921, N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011,
         N1012, N1013, N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021,
         N1022, N1023, N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1031,
         N1032, N1033, N1034, N1035, N1036, N1037, N1038, N1039, N1040, N1041,
         N1042, N1043, N1044, N1045, N1046, N1047, N1048, N1049, N1050, N1051,
         N1052, N1053, N1054, N1055, N1056, N1057, N1058, N1059, N1060, N1061,
         N1062, N1063, N1064, N1065, N1066, N1067, N1068, N1069, N1070, N1071,
         N1072, N1073, N1074, N1075, N1076, N1077, N1078, N1079, N1080, N1081,
         N1082, N1083, N1084, N1085, N1086, N1087, N1088, N1089, N1090, N1091,
         N1092, N1093, N1094, N1095, N1096, N1097, N1098, N1099, N11000, N1101,
         N1102, N1103, N1104, N1105, N1106, N1107, N1108, N1109, N1110, N1111,
         N1112, N1113, N1114, N1115, N1116, N1117, N1118, N1119, N1120, N1121,
         N1122, N1123, N1124, N1125, N1126, N1127, N1128, N1129, N1130, N1131,
         N1132, N1133, N1134, N1135, N1136, N1137, N1138, N1139, N1140, N1141,
         N1142, N1143, N1144, N1145, N1146, N1147, N1148, N1149, N1150, N1151,
         N1152, N1153, N1154, N1155, N1156, N1157, N1158, N1159, N1160, N1161,
         N1162, N1163, N1164, N1165, N1166, N1167, N1168, N1169, N1170, N1171,
         N1172, N1173, N1174, N1175, N1176, N1177, N1178, N1179, N1180, N1181,
         N1182, N1183, N1184, N1185, N1186, N1187, N1188, N1189, N1190, N1191,
         N1192;
  wire   [4:2] CODE_TYPE;
  wire   [2:0] OPER3_R3;
  wire   [3:0] STATE;
  wire   [3:0] NEXT_STATE;
  wire   [15:0] REG_A;
  wire   [15:0] REG_B;
  wire   [12:8] REG_C;

  DFFRX4TF \reg_A_reg[0]  ( .D(N497), .CK(CLK), .RN(RST_N), .Q(REG_A[0]), .QN(
        N213) );
  DFFRX2TF \id_ir_reg[11]  ( .D(N532), .CK(CLK), .RN(RST_N), .Q(N210), .QN(
        N569) );
  DFFRX2TF \gr_reg[3][12]  ( .D(N932), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTB[12]), .QN(N632) );
  DFFRX2TF \gr_reg[1][6]  ( .D(N986), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[6]), 
        .QN(N670) );
  DFFRX2TF \gr_reg[1][5]  ( .D(N987), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[5]), 
        .QN(N671) );
  DFFRX2TF \gr_reg[3][4]  ( .D(N972), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[4]), 
        .QN(N640) );
  DFFRX2TF \gr_reg[3][6]  ( .D(N970), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[6]), 
        .QN(N638) );
  DFFRX2TF \gr_reg[3][5]  ( .D(N971), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[5]), 
        .QN(N639) );
  DFFRX2TF \gr_reg[1][4]  ( .D(N988), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[4]), 
        .QN(N672) );
  DFFRX2TF \gr_reg[3][11]  ( .D(N933), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTB[11]), .QN(N633) );
  DFFRX2TF \gr_reg[3][0]  ( .D(N976), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[0]), 
        .QN(N644) );
  DFFRX2TF \gr_reg[3][15]  ( .D(N929), .CK(CLK), .RN(RST_N), .Q(N242), .QN(
        N629) );
  DFFRX2TF \gr_reg[3][1]  ( .D(N975), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[1]), 
        .QN(N643) );
  DFFRX2TF \gr_reg[3][14]  ( .D(N930), .CK(CLK), .RN(RST_N), .Q(N241), .QN(
        N630) );
  DFFRX2TF \gr_reg[3][10]  ( .D(N934), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTB[10]), .QN(N634) );
  DFFRX2TF \gr_reg[3][9]  ( .D(N935), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[9]), 
        .QN(N635) );
  DFFRX2TF \gr_reg[3][13]  ( .D(N931), .CK(CLK), .RN(RST_N), .Q(N240), .QN(
        N631) );
  DFFRX2TF \gr_reg[3][2]  ( .D(N974), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[2]), 
        .QN(N642) );
  DFFRX2TF \gr_reg[3][8]  ( .D(N936), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[8]), 
        .QN(N636) );
  DFFRX2TF zf_reg ( .D(N434), .CK(CLK), .RN(RST_N), .Q(ZF), .QN(N239) );
  DFFSX2TF \pc_reg[6]  ( .D(N804), .CK(CLK), .SN(RST_N), .Q(N238), .QN(
        I_ADDR[7]) );
  DFFRX2TF \id_ir_reg[8]  ( .D(N535), .CK(CLK), .RN(RST_N), .Q(N236), .QN(N572) );
  DFFSX2TF \pc_reg[4]  ( .D(N809), .CK(CLK), .SN(RST_N), .Q(N235), .QN(
        I_ADDR[5]) );
  DFFSX2TF \pc_reg[1]  ( .D(N812), .CK(CLK), .SN(RST_N), .Q(N234), .QN(
        I_ADDR[2]) );
  DFFRX2TF \reg_A_reg[6]  ( .D(N448), .CK(CLK), .RN(RST_N), .Q(REG_A[6]), .QN(
        N233) );
  DFFRX2TF \reg_A_reg[8]  ( .D(N456), .CK(CLK), .RN(RST_N), .Q(REG_A[8]), .QN(
        N232) );
  DFFRX2TF \reg_A_reg[4]  ( .D(N452), .CK(CLK), .RN(RST_N), .Q(REG_A[4]), .QN(
        N228) );
  DFFRX2TF \gr_reg[3][7]  ( .D(N969), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[7]), 
        .QN(N637) );
  DFFRX2TF \id_ir_reg[4]  ( .D(N523), .CK(CLK), .RN(RST_N), .Q(N227), .QN(N401) );
  DFFRX2TF \id_ir_reg[0]  ( .D(N527), .CK(CLK), .RN(RST_N), .Q(OPER3_R3[0]), 
        .QN(N226) );
  DFFRX2TF \id_ir_reg[10]  ( .D(N533), .CK(CLK), .RN(RST_N), .Q(\OPER1_R1[2] ), 
        .QN(N225) );
  DFFSX2TF \pc_reg[0]  ( .D(N860), .CK(CLK), .SN(RST_N), .Q(N224), .QN(
        I_ADDR[1]) );
  DFFRX2TF \state_reg[3]  ( .D(NEXT_STATE[3]), .CK(CLK), .RN(RST_N), .Q(
        STATE[3]), .QN(N223) );
  DFFRX2TF \reg_A_reg[11]  ( .D(N5070), .CK(CLK), .RN(RST_N), .Q(REG_A[11]), 
        .QN(N222) );
  DFFRX2TF \reg_A_reg[15]  ( .D(N492), .CK(CLK), .RN(RST_N), .Q(REG_A[15]), 
        .QN(N220) );
  DFFRX2TF \id_ir_reg[14]  ( .D(N529), .CK(CLK), .RN(RST_N), .Q(CODE_TYPE[3]), 
        .QN(N219) );
  DFFRX2TF \reg_A_reg[12]  ( .D(N502), .CK(CLK), .RN(RST_N), .Q(REG_A[12]), 
        .QN(N218) );
  DFFRX2TF \reg_A_reg[13]  ( .D(N465), .CK(CLK), .RN(RST_N), .Q(REG_A[13]), 
        .QN(N217) );
  DFFRX2TF \reg_A_reg[2]  ( .D(N461), .CK(CLK), .RN(RST_N), .Q(REG_A[2]), .QN(
        N216) );
  DFFRX2TF \reg_A_reg[7]  ( .D(N5110), .CK(CLK), .RN(RST_N), .Q(REG_A[7]), 
        .QN(N215) );
  DFFRX2TF \reg_A_reg[10]  ( .D(N4740), .CK(CLK), .RN(RST_N), .Q(REG_A[10]), 
        .QN(N214) );
  DFFRX2TF \reg_A_reg[9]  ( .D(N469), .CK(CLK), .RN(RST_N), .Q(REG_A[9]), .QN(
        N212) );
  DFFRX2TF \reg_A_reg[3]  ( .D(N4790), .CK(CLK), .RN(RST_N), .Q(REG_A[3]), 
        .QN(N211) );
  DFFRX2TF \reg_B_reg[3]  ( .D(N4780), .CK(CLK), .RN(RST_N), .Q(REG_B[3]), 
        .QN(N230) );
  DFFRX2TF \id_ir_reg[1]  ( .D(N526), .CK(CLK), .RN(RST_N), .Q(OPER3_R3[1]), 
        .QN(N209) );
  DFFSX2TF \pc_reg[2]  ( .D(N811), .CK(CLK), .SN(RST_N), .Q(N208), .QN(
        I_ADDR[3]) );
  DFFRX2TF \state_reg[1]  ( .D(NEXT_STATE[1]), .CK(CLK), .RN(RST_N), .Q(
        STATE[1]), .QN(N207) );
  DFFRX2TF \id_ir_reg[15]  ( .D(N528), .CK(CLK), .RN(RST_N), .Q(CODE_TYPE[4]), 
        .QN(N206) );
  DFFRX2TF \id_ir_reg[13]  ( .D(N530), .CK(CLK), .RN(RST_N), .Q(CODE_TYPE[2]), 
        .QN(N205) );
  DFFRX2TF \id_ir_reg[2]  ( .D(N525), .CK(CLK), .RN(RST_N), .Q(OPER3_R3[2]), 
        .QN(N204) );
  DFFRX2TF \state_reg[2]  ( .D(NEXT_STATE[2]), .CK(CLK), .RN(RST_N), .Q(N203), 
        .QN(N554) );
  DFFRX2TF \reg_A_reg[14]  ( .D(N4830), .CK(CLK), .RN(RST_N), .Q(REG_A[14]), 
        .QN(N202) );
  DFFRX2TF \reg_A_reg[5]  ( .D(N444), .CK(CLK), .RN(RST_N), .Q(REG_A[5]), .QN(
        N201) );
  DFFRX2TF \reg_A_reg[1]  ( .D(N488), .CK(CLK), .RN(RST_N), .Q(REG_A[1]), .QN(
        N200) );
  TLATXLTF cf_buf_reg ( .G(N588), .D(N589), .Q(CF_BUF) );
  TLATXLTF \nxt_reg[0]  ( .G(N166), .D(N167), .Q(NXT[0]) );
  TLATXLTF \nxt_reg[1]  ( .G(N166), .D(N168), .Q(NXT[1]) );
  DFFRX2TF \gr_reg[4][9]  ( .D(N927), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[9]), 
        .QN(N619) );
  DFFRX2TF \gr_reg[4][7]  ( .D(N961), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[7]), 
        .QN(N621) );
  DFFRX2TF \gr_reg[4][8]  ( .D(N928), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[8]), 
        .QN(N620) );
  DFFRX2TF \gr_reg[4][6]  ( .D(N962), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[6]), 
        .QN(N622) );
  DFFRX2TF \gr_reg[4][5]  ( .D(N963), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[5]), 
        .QN(N623) );
  DFFRX2TF \gr_reg[4][1]  ( .D(N967), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[1]), 
        .QN(N627) );
  DFFRX2TF \gr_reg[4][3]  ( .D(N965), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[3]), 
        .QN(N625) );
  DFFRX2TF \gr_reg[4][2]  ( .D(N966), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[2]), 
        .QN(N626) );
  DFFRX2TF \gr_reg[4][4]  ( .D(N964), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[4]), 
        .QN(N624) );
  DFFRX2TF \gr_reg[4][0]  ( .D(N968), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[0]), 
        .QN(N628) );
  DFFSX2TF \pc_reg[5]  ( .D(N808), .CK(CLK), .SN(RST_N), .QN(I_ADDR[6]) );
  DFFSX2TF \pc_reg[7]  ( .D(N859), .CK(CLK), .SN(RST_N), .QN(I_ADDR[8]) );
  DFFSX2TF \pc_reg[3]  ( .D(N810), .CK(CLK), .SN(RST_N), .QN(I_ADDR[4]) );
  DFFRX2TF \gr_reg[1][0]  ( .D(N992), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[0]), 
        .QN(N676) );
  DFFRX2TF \gr_reg[1][1]  ( .D(N991), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[1]), 
        .QN(N675) );
  DFFRX2TF \gr_reg[2][11]  ( .D(N941), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTA[11]), .QN(N649) );
  DFFRX2TF \reg_B_reg[14]  ( .D(N437), .CK(CLK), .RN(RST_N), .Q(REG_B[14]), 
        .QN(N415) );
  DFFRX2TF \reg_B_reg[15]  ( .D(N436), .CK(CLK), .RN(RST_N), .Q(REG_B[15]), 
        .QN(N412) );
  DFFRX2TF \gr_reg[2][12]  ( .D(N940), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTA[12]), .QN(N648) );
  DFFRX2TF \gr_reg[2][8]  ( .D(N944), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[8]), 
        .QN(N652) );
  DFFRX2TF \gr_reg[2][10]  ( .D(N942), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTA[10]), .QN(N650) );
  DFFRX2TF \gr_reg[2][9]  ( .D(N943), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[9]), 
        .QN(N651) );
  DFFRX2TF \reg_B_reg[11]  ( .D(N5060), .CK(CLK), .RN(RST_N), .Q(REG_B[11]), 
        .QN(N409) );
  DFFRX2TF \reg_B_reg[12]  ( .D(N501), .CK(CLK), .RN(RST_N), .Q(REG_B[12]), 
        .QN(N411) );
  DFFRX2TF \reg_B_reg[10]  ( .D(N4730), .CK(CLK), .RN(RST_N), .Q(REG_B[10]), 
        .QN(N408) );
  DFFRX2TF \reg_B_reg[13]  ( .D(N439), .CK(CLK), .RN(RST_N), .Q(REG_B[13]), 
        .QN(N413) );
  DFFRX2TF \reg_B_reg[9]  ( .D(N438), .CK(CLK), .RN(RST_N), .Q(REG_B[9]), .QN(
        N418) );
  DFFRX2TF \gr_reg[2][3]  ( .D(N981), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[3]), 
        .QN(N657) );
  DFFRX2TF \gr_reg[2][5]  ( .D(N979), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[5]), 
        .QN(N655) );
  DFFRX2TF \gr_reg[1][2]  ( .D(N990), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[2]), 
        .QN(N674) );
  DFFRX2TF \gr_reg[1][3]  ( .D(N989), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[3]), 
        .QN(N673) );
  DFFRX2TF \gr_reg[2][1]  ( .D(N983), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[1]), 
        .QN(N659) );
  DFFRX2TF \gr_reg[2][6]  ( .D(N978), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[6]), 
        .QN(N654) );
  DFFRX2TF \gr_reg[2][2]  ( .D(N982), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[2]), 
        .QN(N658) );
  DFFRX2TF \gr_reg[2][7]  ( .D(N977), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[7]), 
        .QN(N653) );
  DFFRX2TF \gr_reg[2][4]  ( .D(N980), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[4]), 
        .QN(N656) );
  DFFRX2TF \reg_B_reg[7]  ( .D(N5140), .CK(CLK), .RN(RST_N), .Q(REG_B[7]), 
        .QN(N405) );
  DFFRX2TF \reg_B_reg[5]  ( .D(N443), .CK(CLK), .RN(RST_N), .Q(REG_B[5]), .QN(
        N424) );
  DFFRX2TF \reg_B_reg[6]  ( .D(N442), .CK(CLK), .RN(RST_N), .Q(REG_B[6]), .QN(
        N406) );
  DFFRX2TF \reg_B_reg[8]  ( .D(N440), .CK(CLK), .RN(RST_N), .Q(REG_B[8]), .QN(
        N420) );
  DFFRX2TF \gr_reg[2][0]  ( .D(N984), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[0]), 
        .QN(N660) );
  DFFRX2TF \gr_reg[3][3]  ( .D(N973), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[3]), 
        .QN(N641) );
  DFFRX2TF \state_reg[0]  ( .D(NEXT_STATE[0]), .CK(CLK), .RN(RST_N), .Q(
        STATE[0]), .QN(N231) );
  DFFRX2TF \reg_B_reg[4]  ( .D(N441), .CK(CLK), .RN(RST_N), .Q(REG_B[4]), .QN(
        N423) );
  CMPR32X2TF \sub_x_285_4/U9  ( .A(N420), .B(REG_A[8]), .C(SUB_X_285_4_N9), 
        .CO(SUB_X_285_4_N8), .S(N512) );
  CMPR32X2TF \sub_x_285_4/U6  ( .A(N409), .B(REG_A[11]), .C(SUB_X_285_4_N6), 
        .CO(SUB_X_285_4_N5), .S(N515) );
  CMPR32X2TF \sub_x_285_4/U10  ( .A(N405), .B(REG_A[7]), .C(SUB_X_285_4_N10), 
        .CO(SUB_X_285_4_N9), .S(N511) );
  CMPR32X2TF \sub_x_285_4/U12  ( .A(N424), .B(REG_A[5]), .C(SUB_X_285_4_N12), 
        .CO(SUB_X_285_4_N11), .S(N509) );
  CMPR32X2TF \sub_x_285_4/U11  ( .A(N406), .B(REG_A[6]), .C(SUB_X_285_4_N11), 
        .CO(SUB_X_285_4_N10), .S(N510) );
  CMPR32X2TF \sub_x_285_4/U5  ( .A(N411), .B(REG_A[12]), .C(SUB_X_285_4_N5), 
        .CO(SUB_X_285_4_N4), .S(N516) );
  CMPR32X2TF \sub_x_285_4/U16  ( .A(N193), .B(REG_A[1]), .C(SUB_X_285_4_N16), 
        .CO(SUB_X_285_4_N15), .S(N505) );
  CMPR32X2TF \sub_x_285_4/U4  ( .A(N413), .B(REG_A[13]), .C(SUB_X_285_4_N4), 
        .CO(SUB_X_285_4_N3), .S(N517) );
  CMPR32X2TF \sub_x_285_4/U3  ( .A(N415), .B(REG_A[14]), .C(SUB_X_285_4_N3), 
        .CO(SUB_X_285_4_N2), .S(N518) );
  CMPR32X2TF \add_x_285_3/U5  ( .A(REG_A[12]), .B(REG_B[12]), .C(
        ADD_X_285_3_N5), .CO(ADD_X_285_3_N4), .S(N482) );
  CMPR32X2TF \add_x_285_3/U6  ( .A(REG_A[11]), .B(REG_B[11]), .C(
        ADD_X_285_3_N6), .CO(ADD_X_285_3_N5), .S(N481) );
  CMPR32X2TF \add_x_285_3/U7  ( .A(REG_A[10]), .B(REG_B[10]), .C(
        ADD_X_285_3_N7), .CO(ADD_X_285_3_N6), .S(N480) );
  CMPR32X2TF \add_x_285_3/U3  ( .A(REG_A[14]), .B(REG_B[14]), .C(
        ADD_X_285_3_N3), .CO(ADD_X_285_3_N2), .S(N484) );
  CMPR32X2TF \add_x_285_3/U16  ( .A(REG_A[1]), .B(REG_B[1]), .C(
        ADD_X_285_3_N16), .CO(ADD_X_285_3_N15), .S(N471) );
  CMPR32X2TF \add_x_285_3/U15  ( .A(REG_A[2]), .B(N142), .C(ADD_X_285_3_N15), 
        .CO(ADD_X_285_3_N14), .S(N472) );
  CMPR32X2TF \add_x_285_3/U14  ( .A(REG_A[3]), .B(REG_B[3]), .C(
        ADD_X_285_3_N14), .CO(ADD_X_285_3_N13), .S(N473) );
  CMPR32X2TF \add_x_285_3/U13  ( .A(REG_A[4]), .B(REG_B[4]), .C(
        ADD_X_285_3_N13), .CO(ADD_X_285_3_N12), .S(N474) );
  CMPR32X2TF \add_x_285_3/U12  ( .A(REG_A[5]), .B(REG_B[5]), .C(
        ADD_X_285_3_N12), .CO(ADD_X_285_3_N11), .S(N475) );
  CMPR32X2TF \add_x_285_3/U11  ( .A(REG_A[6]), .B(REG_B[6]), .C(
        ADD_X_285_3_N11), .CO(ADD_X_285_3_N10), .S(N476) );
  CMPR32X2TF \add_x_285_3/U10  ( .A(REG_A[7]), .B(REG_B[7]), .C(
        ADD_X_285_3_N10), .CO(ADD_X_285_3_N9), .S(N477) );
  CMPR32X2TF \add_x_285_3/U9  ( .A(REG_A[8]), .B(REG_B[8]), .C(ADD_X_285_3_N9), 
        .CO(ADD_X_285_3_N8), .S(N478) );
  CMPR32X2TF \add_x_285_3/U8  ( .A(REG_A[9]), .B(REG_B[9]), .C(ADD_X_285_3_N8), 
        .CO(ADD_X_285_3_N7), .S(N479) );
  CMPR32X2TF \add_x_285_3/U4  ( .A(REG_A[13]), .B(REG_B[13]), .C(
        ADD_X_285_3_N4), .CO(ADD_X_285_3_N3), .S(N483) );
  DFFNSRX2TF lowest_bit_reg ( .D(N1002), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        I_ADDR[0]), .QN(N221) );
  DFFNSRXLTF \reg_C_reg[13]  ( .D(N468), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N421) );
  DFFNSRXLTF \reg_C_reg[14]  ( .D(N4860), .CKN(CLK), .SN(1'b1), .RN(1'b1), 
        .QN(N416) );
  DFFNSRXLTF \reg_C_reg[15]  ( .D(N495), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N414) );
  DFFNSRXLTF is_i_addr_reg ( .D(N110), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        IS_I_ADDR) );
  DFFNSRXLTF dw_reg ( .D(N616), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(D_WE) );
  DFFNSRXLTF \reg_C_reg[9]  ( .D(N4720), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        REG_C[9]) );
  DFFNSRXLTF \reg_C_reg[11]  ( .D(N5100), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        REG_C[11]) );
  DFFNSRXLTF \reg_C_reg[12]  ( .D(N5050), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        REG_C[12]) );
  DFFNSRXLTF \reg_C_reg[8]  ( .D(N459), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        REG_C[8]) );
  DFFNSRXLTF \reg_C_reg[10]  ( .D(N4770), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        REG_C[10]) );
  DFFRX4TF \reg_B_reg[0]  ( .D(N496), .CK(CLK), .RN(RST_N), .Q(REG_B[0]), .QN(
        N1129) );
  DFFRX1TF \smdr_reg[9]  ( .D(N4700), .CK(CLK), .RN(RST_N), .QN(N601) );
  DFFRX1TF \smdr_reg[8]  ( .D(N457), .CK(CLK), .RN(RST_N), .QN(N602) );
  DFFRX1TF \smdr_reg[6]  ( .D(N449), .CK(CLK), .RN(RST_N), .QN(N604) );
  DFFRX1TF \smdr_reg[5]  ( .D(N445), .CK(CLK), .RN(RST_N), .QN(N605) );
  DFFRX1TF \smdr_reg[4]  ( .D(N453), .CK(CLK), .RN(RST_N), .QN(N606) );
  DFFRX1TF \smdr_reg[2]  ( .D(N462), .CK(CLK), .RN(RST_N), .QN(N608) );
  DFFRX1TF \smdr_reg[1]  ( .D(N489), .CK(CLK), .RN(RST_N), .QN(N609) );
  DFFRX1TF \smdr_reg[15]  ( .D(N493), .CK(CLK), .RN(RST_N), .QN(N595) );
  DFFRX1TF \smdr_reg[14]  ( .D(N4840), .CK(CLK), .RN(RST_N), .QN(N596) );
  DFFRX1TF \smdr_reg[13]  ( .D(N466), .CK(CLK), .RN(RST_N), .QN(N597) );
  DFFRX1TF \smdr_reg[12]  ( .D(N503), .CK(CLK), .RN(RST_N), .QN(N598) );
  DFFRX1TF \smdr_reg[11]  ( .D(N5080), .CK(CLK), .RN(RST_N), .QN(N599) );
  DFFRX1TF \smdr_reg[10]  ( .D(N4750), .CK(CLK), .RN(RST_N), .QN(N600) );
  DFFRX1TF \smdr_reg[7]  ( .D(N433), .CK(CLK), .RN(RST_N), .QN(N603) );
  DFFRX1TF \smdr_reg[3]  ( .D(N4800), .CK(CLK), .RN(RST_N), .QN(N607) );
  DFFRX1TF \smdr_reg[0]  ( .D(N498), .CK(CLK), .RN(RST_N), .QN(N610) );
  DFFRX1TF nf_reg ( .D(N435), .CK(CLK), .RN(RST_N), .QN(N237) );
  DFFRX1TF \id_ir_reg[7]  ( .D(N520), .CK(CLK), .RN(RST_N), .QN(N404) );
  DFFRX1TF \id_ir_reg[3]  ( .D(N524), .CK(CLK), .RN(RST_N), .QN(N400) );
  DFFRX1TF \id_ir_reg[6]  ( .D(N521), .CK(CLK), .RN(RST_N), .QN(N403) );
  DFFRX1TF \id_ir_reg[5]  ( .D(N522), .CK(CLK), .RN(RST_N), .QN(N402) );
  DFFRX1TF \gr_reg[0][15]  ( .D(N953), .CK(CLK), .RN(RST_N), .QN(N677) );
  DFFRX1TF \gr_reg[0][14]  ( .D(N954), .CK(CLK), .RN(RST_N), .QN(N678) );
  DFFRX1TF \gr_reg[0][13]  ( .D(N955), .CK(CLK), .RN(RST_N), .QN(N679) );
  DFFRX1TF \gr_reg[4][15]  ( .D(N1001), .CK(CLK), .RN(RST_N), .QN(N613) );
  DFFRX1TF \gr_reg[4][14]  ( .D(N922), .CK(CLK), .RN(RST_N), .QN(N614) );
  DFFRX1TF \gr_reg[4][13]  ( .D(N923), .CK(CLK), .RN(RST_N), .QN(N615) );
  DFFRX1TF \gr_reg[2][15]  ( .D(N937), .CK(CLK), .RN(RST_N), .QN(N645) );
  DFFRX1TF \gr_reg[2][14]  ( .D(N938), .CK(CLK), .RN(RST_N), .QN(N646) );
  DFFRX1TF \gr_reg[2][13]  ( .D(N939), .CK(CLK), .RN(RST_N), .QN(N647) );
  DFFRX1TF \gr_reg[1][15]  ( .D(N945), .CK(CLK), .RN(RST_N), .QN(N661) );
  DFFRX1TF \gr_reg[1][14]  ( .D(N946), .CK(CLK), .RN(RST_N), .QN(N662) );
  DFFRX1TF \gr_reg[1][13]  ( .D(N947), .CK(CLK), .RN(RST_N), .QN(N663) );
  DFFRX1TF \gr_reg[0][12]  ( .D(N956), .CK(CLK), .RN(RST_N), .QN(N680) );
  DFFRX1TF \gr_reg[0][11]  ( .D(N957), .CK(CLK), .RN(RST_N), .QN(N681) );
  DFFRX1TF \gr_reg[0][10]  ( .D(N958), .CK(CLK), .RN(RST_N), .QN(N682) );
  DFFRX1TF \gr_reg[0][9]  ( .D(N959), .CK(CLK), .RN(RST_N), .QN(N683) );
  DFFRX1TF \gr_reg[0][8]  ( .D(N960), .CK(CLK), .RN(RST_N), .QN(N684) );
  DFFRX1TF \gr_reg[0][4]  ( .D(N996), .CK(CLK), .RN(RST_N), .QN(N688) );
  DFFRX1TF \gr_reg[0][3]  ( .D(N997), .CK(CLK), .RN(RST_N), .QN(N689) );
  DFFRX1TF \gr_reg[0][2]  ( .D(N998), .CK(CLK), .RN(RST_N), .QN(N690) );
  DFFRX1TF \gr_reg[0][1]  ( .D(N999), .CK(CLK), .RN(RST_N), .QN(N691) );
  DFFRX1TF \gr_reg[0][0]  ( .D(N1000), .CK(CLK), .RN(RST_N), .QN(N692) );
  DFFRX1TF \gr_reg[4][12]  ( .D(N924), .CK(CLK), .RN(RST_N), .QN(N6160) );
  DFFRX1TF \gr_reg[4][11]  ( .D(N925), .CK(CLK), .RN(RST_N), .QN(N617) );
  DFFRX1TF \gr_reg[4][10]  ( .D(N926), .CK(CLK), .RN(RST_N), .QN(N618) );
  DFFRX1TF \gr_reg[0][7]  ( .D(N993), .CK(CLK), .RN(RST_N), .QN(N685) );
  DFFRX1TF \gr_reg[0][6]  ( .D(N994), .CK(CLK), .RN(RST_N), .QN(N686) );
  DFFRX1TF \gr_reg[0][5]  ( .D(N995), .CK(CLK), .RN(RST_N), .QN(N687) );
  DFFRX1TF \gr_reg[1][12]  ( .D(N948), .CK(CLK), .RN(RST_N), .QN(N664) );
  DFFRX1TF \gr_reg[1][11]  ( .D(N949), .CK(CLK), .RN(RST_N), .QN(N665) );
  DFFRX1TF \gr_reg[1][10]  ( .D(N950), .CK(CLK), .RN(RST_N), .QN(N666) );
  DFFRX1TF \gr_reg[1][9]  ( .D(N951), .CK(CLK), .RN(RST_N), .QN(N667) );
  DFFRX1TF \gr_reg[1][8]  ( .D(N952), .CK(CLK), .RN(RST_N), .QN(N668) );
  DFFRX1TF \gr_reg[1][7]  ( .D(N985), .CK(CLK), .RN(RST_N), .QN(N669) );
  DFFRX1TF cf_reg ( .D(N5180), .CK(CLK), .RN(RST_N), .Q(CF) );
  DFFRX1TF \reg_B_reg[2]  ( .D(N460), .CK(CLK), .RN(RST_N), .Q(N43), .QN(N141)
         );
  DFFRX2TF \id_ir_reg[9]  ( .D(N534), .CK(CLK), .RN(RST_N), .Q(N736), .QN(N571) );
  DFFNSRX2TF \reg_C_reg[2]  ( .D(N464), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[3]) );
  DFFNSRX2TF \reg_C_reg[6]  ( .D(N451), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[7]) );
  DFFNSRX2TF \reg_C_reg[4]  ( .D(N455), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[5]) );
  DFFNSRX2TF \reg_C_reg[5]  ( .D(N447), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[6]) );
  DFFNSRX2TF \reg_C_reg[1]  ( .D(N491), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[2]) );
  DFFNSRX2TF \reg_C_reg[3]  ( .D(N4820), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[4]) );
  DFFNSRX1TF \reg_C_reg[0]  ( .D(N500), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[1]) );
  DFFNSRX2TF \reg_C_reg[7]  ( .D(N5130), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[8]) );
  DFFRX2TF \id_ir_reg[12]  ( .D(N531), .CK(CLK), .RN(RST_N), .Q(N250), .QN(N42) );
  DFFRX2TF \reg_B_reg[1]  ( .D(N487), .CK(CLK), .RN(RST_N), .Q(REG_B[1]), .QN(
        N193) );
  AOI21X2TF U3 ( .A0(N483), .A1(N348), .B0(N277), .Y(N397) );
  NAND2X1TF U4 ( .A(N398), .B(N230), .Y(N335) );
  CMPR32X2TF U5 ( .A(N412), .B(REG_A[15]), .C(SUB_X_285_4_N2), .CO(
        SUB_X_285_4_N1), .S(N519) );
  ADDFX2TF U6 ( .A(REG_A[15]), .B(REG_B[15]), .CI(ADD_X_285_3_N2), .CO(N486), 
        .S(N485) );
  OAI21X1TF U7 ( .A0(N381), .A1(N147), .B0(N380), .Y(N500) );
  AO21X1TF U8 ( .A0(N407), .A1(N405), .B0(N143), .Y(N1) );
  OAI222X1TF U9 ( .A0(N795), .A1(N835), .B0(N797), .B1(N837), .C0(N794), .C1(
        N864), .Y(N2) );
  OAI2BB2XLTF U10 ( .B0(N802), .B1(N833), .A0N(N341), .A1N(N332), .Y(N3) );
  AOI211X1TF U11 ( .A0(REG_A[7]), .A1(N1), .B0(N2), .C0(N3), .Y(N4) );
  AOI22X1TF U12 ( .A0(REG_A[7]), .A1(N175), .B0(N252), .B1(N215), .Y(N5) );
  AOI32X1TF U13 ( .A0(N156), .A1(N4), .A2(N5), .B0(N405), .B1(N4), .Y(N6) );
  AO21X1TF U14 ( .A0(N244), .A1(N511), .B0(N6), .Y(N7) );
  AOI21X1TF U15 ( .A0(N348), .A1(N477), .B0(N7), .Y(N385) );
  AOI2BB2X1TF U16 ( .B0(N1173), .B1(IO_DATAINA[10]), .A0N(N372), .A1N(N146), 
        .Y(N8) );
  AOI22X1TF U17 ( .A0(N1171), .A1(REG_C[10]), .B0(N389), .B1(IO_DATAINB[10]), 
        .Y(N9) );
  OAI211X1TF U18 ( .A0(N382), .A1(N149), .B0(N8), .C0(N9), .Y(N4770) );
  AO21X1TF U19 ( .A0(N407), .A1(N423), .B0(N143), .Y(N10) );
  AOI22X1TF U20 ( .A0(N348), .A1(N474), .B0(N865), .B1(N508), .Y(N11) );
  OA22X1TF U21 ( .A0(N837), .A1(N825), .B0(N864), .B1(N824), .Y(N12) );
  OAI211X1TF U22 ( .A0(N833), .A1(N834), .B0(N11), .C0(N12), .Y(N13) );
  CLKINVX1TF U23 ( .A(N341), .Y(N14) );
  CLKINVX1TF U24 ( .A(N854), .Y(N15) );
  OAI22X1TF U25 ( .A0(N832), .A1(N14), .B0(N846), .B1(N15), .Y(N16) );
  AOI211X1TF U26 ( .A0(REG_A[4]), .A1(N10), .B0(N13), .C0(N16), .Y(N17) );
  AOI22X1TF U27 ( .A0(REG_A[4]), .A1(N175), .B0(N407), .B1(N228), .Y(N18) );
  AOI32X1TF U28 ( .A0(N157), .A1(N17), .A2(N18), .B0(N423), .B1(N17), .Y(N361)
         );
  AOI2BB2X1TF U29 ( .B0(N1173), .B1(IO_DATAINA[11]), .A0N(N382), .A1N(N146), 
        .Y(N19) );
  AOI22X1TF U30 ( .A0(N1171), .A1(REG_C[11]), .B0(N246), .B1(IO_DATAINB[11]), 
        .Y(N20) );
  OAI211X1TF U31 ( .A0(N383), .A1(N149), .B0(N19), .C0(N20), .Y(N5100) );
  AOI22X1TF U32 ( .A0(REG_A[6]), .A1(N175), .B0(N252), .B1(N233), .Y(N21) );
  AOI21X1TF U33 ( .A0(N157), .A1(N21), .B0(N406), .Y(N22) );
  AOI21X1TF U34 ( .A0(N251), .A1(N406), .B0(N143), .Y(N23) );
  OAI22X1TF U35 ( .A0(N872), .A1(N864), .B0(N742), .B1(N784), .Y(N24) );
  OAI2BB2XLTF U36 ( .B0(N835), .B1(N779), .A0N(N782), .A1N(N840), .Y(N25) );
  AOI211X1TF U37 ( .A0(N865), .A1(N510), .B0(N24), .C0(N25), .Y(N26) );
  OAI21X1TF U38 ( .A0(N233), .A1(N23), .B0(N26), .Y(N27) );
  AOI211X1TF U39 ( .A0(N348), .A1(N476), .B0(N22), .C0(N27), .Y(N28) );
  OAI21X1TF U40 ( .A0(N831), .A1(N863), .B0(N28), .Y(N387) );
  AOI2BB2X1TF U41 ( .B0(N1173), .B1(IO_DATAINA[12]), .A0N(N383), .A1N(N146), 
        .Y(N29) );
  AOI22X1TF U42 ( .A0(N1171), .A1(REG_C[12]), .B0(N246), .B1(IO_DATAINB[12]), 
        .Y(N30) );
  OAI211X1TF U43 ( .A0(N396), .A1(N149), .B0(N29), .C0(N30), .Y(N5050) );
  AOI2BB1X1TF U44 ( .A0N(N145), .A1N(N835), .B0(N5090), .Y(N320) );
  OAI21X1TF U45 ( .A0(N774), .A1(N212), .B0(N745), .Y(N31) );
  NOR3X1TF U46 ( .A(N743), .B(N744), .C(N31), .Y(N779) );
  AOI2BB2X1TF U47 ( .B0(N227), .B1(N1021), .A0N(N1025), .A1N(N1020), .Y(N163)
         );
  OA21XLTF U48 ( .A0(N708), .A1(I_ADDR[4]), .B0(N709), .Y(N32) );
  AOI222XLTF U49 ( .A0(I_ADDR[4]), .A1(N714), .B0(N721), .B1(D_ADDR[4]), .C0(
        N712), .C1(N32), .Y(N810) );
  CLKINVX1TF U50 ( .A(N244), .Y(N33) );
  OAI22X1TF U51 ( .A0(SUB_X_285_4_N1), .A1(N33), .B0(N34), .B1(N538), .Y(N589)
         );
  CLKINVX1TF U52 ( .A(N486), .Y(N34) );
  NAND2BX1TF U53 ( .AN(N878), .B(N1004), .Y(N35) );
  OAI211X1TF U54 ( .A0(N1006), .A1(N419), .B0(N1005), .C0(N35), .Y(N1016) );
  OA21XLTF U55 ( .A0(N713), .A1(I_ADDR[6]), .B0(N718), .Y(N36) );
  AOI222XLTF U56 ( .A0(I_ADDR[6]), .A1(N714), .B0(N721), .B1(D_ADDR[6]), .C0(
        N712), .C1(N36), .Y(N808) );
  NOR4XLTF U57 ( .A(N1186), .B(N355), .C(N356), .D(N361), .Y(N37) );
  NAND4X1TF U58 ( .A(N37), .B(N385), .C(N390), .D(N392), .Y(N38) );
  NOR4XLTF U59 ( .A(N368), .B(N387), .C(N363), .D(N38), .Y(N39) );
  AND4X1TF U60 ( .A(N39), .B(N372), .C(N382), .D(N383), .Y(N40) );
  NAND4X1TF U61 ( .A(N40), .B(N396), .C(N397), .D(N395), .Y(N41) );
  OAI2BB2XLTF U62 ( .B0(N376), .B1(N41), .A0N(N1186), .A1N(ZF), .Y(N434) );
  OR2X2TF U63 ( .A(N193), .B(REG_B[0]), .Y(N44) );
  OR3X1TF U64 ( .A(N1006), .B(N879), .C(N42), .Y(N869) );
  CLKBUFX2TF U65 ( .A(N1179), .Y(N53) );
  INVX1TF U85 ( .A(N846), .Y(N852) );
  CLKINVX4TF U86 ( .A(N407), .Y(N139) );
  CLKINVX2TF U87 ( .A(N555), .Y(N264) );
  OR3X1TF U88 ( .A(N741), .B(N877), .C(N875), .Y(N1159) );
  INVX4TF U89 ( .A(N142), .Y(N140) );
  NAND2XLTF U90 ( .A(N419), .B(CODE_TYPE[3]), .Y(N880) );
  INVX2TF U91 ( .A(N250), .Y(N158) );
  XOR2X1TF U92 ( .A(N396), .B(N382), .Y(N374) );
  AO22X1TF U93 ( .A0(N1023), .A1(N1022), .B0(N401), .B1(N1021), .Y(N1166) );
  OAI22X1TF U94 ( .A0(N225), .A1(N1025), .B0(N1024), .B1(N403), .Y(N1165) );
  OAI31XLTF U95 ( .A0(IO_STATUS[0]), .A1(IO_STATUS[1]), .A2(N732), .B0(N731), 
        .Y(NEXT_STATE[1]) );
  NAND4X2TF U96 ( .A(N226), .B(N209), .C(N204), .D(N887), .Y(N1175) );
  INVX2TF U97 ( .A(N887), .Y(N888) );
  NAND2X1TF U98 ( .A(N230), .B(N866), .Y(N868) );
  OAI211XLTF U99 ( .A0(N1034), .A1(N1006), .B0(N552), .C0(N551), .Y(N553) );
  NAND2XLTF U100 ( .A(N422), .B(REG_A[5]), .Y(N763) );
  INVX2TF U101 ( .A(N144), .Y(N422) );
  INVX2TF U102 ( .A(N735), .Y(N730) );
  CMPR22X2TF U103 ( .A(REG_B[0]), .B(REG_A[0]), .CO(ADD_X_285_3_N16), .S(N470)
         );
  OAI222X1TF U104 ( .A0(N149), .A1(N373), .B0(N147), .B1(N395), .C0(N414), 
        .C1(N243), .Y(N495) );
  AOI22X1TF U105 ( .A0(N568), .A1(N576), .B0(N641), .B1(N567), .Y(N973) );
  AOI22X1TF U106 ( .A0(N563), .A1(N576), .B0(N673), .B1(N562), .Y(N989) );
  AOI22X1TF U107 ( .A0(N565), .A1(N574), .B0(N659), .B1(N564), .Y(N983) );
  AOI22X1TF U108 ( .A0(N565), .A1(N573), .B0(N660), .B1(N564), .Y(N984) );
  AOI21X1TF U109 ( .A0(N480), .A1(N245), .B0(N313), .Y(N382) );
  AOI22X1TF U110 ( .A0(N693), .A1(N698), .B0(N632), .B1(N611), .Y(N932) );
  AOI22X1TF U111 ( .A0(N568), .A1(N577), .B0(N640), .B1(N567), .Y(N972) );
  AOI22X1TF U112 ( .A0(N565), .A1(N577), .B0(N656), .B1(N564), .Y(N980) );
  AOI22X1TF U113 ( .A0(N693), .A1(N697), .B0(N633), .B1(N611), .Y(N933) );
  AOI22X1TF U114 ( .A0(N593), .A1(N697), .B0(N649), .B1(N592), .Y(N941) );
  AOI22X1TF U115 ( .A0(N568), .A1(N573), .B0(N644), .B1(N567), .Y(N976) );
  AOI22X1TF U116 ( .A0(N563), .A1(N574), .B0(N675), .B1(N562), .Y(N991) );
  AOI22X1TF U117 ( .A0(N563), .A1(N573), .B0(N676), .B1(N562), .Y(N992) );
  AOI22X1TF U118 ( .A0(N568), .A1(N574), .B0(N643), .B1(N567), .Y(N975) );
  AOI22X1TF U119 ( .A0(N591), .A1(N695), .B0(N667), .B1(N590), .Y(N951) );
  AOI22X1TF U120 ( .A0(N693), .A1(N696), .B0(N634), .B1(N611), .Y(N934) );
  AOI22X1TF U121 ( .A0(N693), .A1(N695), .B0(N635), .B1(N611), .Y(N935) );
  AOI22X1TF U122 ( .A0(N591), .A1(N696), .B0(N666), .B1(N590), .Y(N950) );
  AOI22X1TF U123 ( .A0(N591), .A1(N698), .B0(N664), .B1(N590), .Y(N948) );
  AOI22X1TF U124 ( .A0(N593), .A1(N695), .B0(N651), .B1(N592), .Y(N943) );
  AOI22X1TF U125 ( .A0(N593), .A1(N696), .B0(N650), .B1(N592), .Y(N942) );
  AOI22X1TF U126 ( .A0(N593), .A1(N698), .B0(N648), .B1(N592), .Y(N940) );
  NOR4XLTF U127 ( .A(N822), .B(N344), .C(N823), .D(N343), .Y(N345) );
  OAI22X1TF U128 ( .A0(N683), .A1(N189), .B0(N651), .B1(N186), .Y(N1077) );
  OAI22X1TF U129 ( .A0(N677), .A1(N189), .B0(N645), .B1(N186), .Y(N1125) );
  OAI22X1TF U130 ( .A0(N169), .A1(N601), .B0(N667), .B1(N183), .Y(N1078) );
  OAI22X1TF U131 ( .A0(N679), .A1(N190), .B0(N647), .B1(N187), .Y(N1071) );
  OAI22X1TF U132 ( .A0(N684), .A1(N189), .B0(N652), .B1(N186), .Y(N1053) );
  OAI22X1TF U133 ( .A0(N678), .A1(N190), .B0(N646), .B1(N187), .Y(N1105) );
  OAI22X1TF U134 ( .A0(N170), .A1(N602), .B0(N668), .B1(N183), .Y(N1054) );
  OAI22X1TF U135 ( .A0(N680), .A1(N190), .B0(N648), .B1(N187), .Y(N1148) );
  OAI22X1TF U136 ( .A0(N682), .A1(N190), .B0(N650), .B1(N187), .Y(N1087) );
  OAI22X1TF U137 ( .A0(N631), .A1(N191), .B0(N663), .B1(N1177), .Y(N903) );
  OAI22X1TF U138 ( .A0(N681), .A1(N190), .B0(N649), .B1(N187), .Y(N1160) );
  OAI22X1TF U139 ( .A0(N692), .A1(N190), .B0(N660), .B1(N187), .Y(N1137) );
  NAND3XLTF U140 ( .A(N539), .B(N845), .C(N538), .Y(N588) );
  AO22X1TF U141 ( .A0(N227), .A1(N1019), .B0(N1018), .B1(N1022), .Y(N1164) );
  OAI22X1TF U142 ( .A0(N685), .A1(N190), .B0(N653), .B1(N187), .Y(N737) );
  OAI22X1TF U143 ( .A0(N691), .A1(N189), .B0(N659), .B1(N186), .Y(N1115) );
  OAI22X1TF U144 ( .A0(N689), .A1(N190), .B0(N657), .B1(N187), .Y(N1097) );
  OAI22X1TF U145 ( .A0(N170), .A1(N608), .B0(N674), .B1(N183), .Y(N1064) );
  OAI22X1TF U146 ( .A0(N629), .A1(N191), .B0(N661), .B1(N1177), .Y(N891) );
  OAI22X1TF U147 ( .A0(N690), .A1(N189), .B0(N658), .B1(N186), .Y(N1063) );
  OAI22X1TF U148 ( .A0(N687), .A1(N189), .B0(N655), .B1(N186), .Y(N1029) );
  OAI22X1TF U149 ( .A0(N169), .A1(N606), .B0(N672), .B1(N183), .Y(N1047) );
  OAI22X1TF U150 ( .A0(N170), .A1(N605), .B0(N671), .B1(N183), .Y(N1030) );
  OAI22X1TF U151 ( .A0(N688), .A1(N189), .B0(N656), .B1(N186), .Y(N1046) );
  OAI22X1TF U152 ( .A0(N630), .A1(N191), .B0(N662), .B1(N1177), .Y(N895) );
  OAI22X1TF U153 ( .A0(N614), .A1(N1660), .B0(N646), .B1(N1180), .Y(N894) );
  OAI22X1TF U154 ( .A0(N1680), .A1(N604), .B0(N670), .B1(N183), .Y(N1041) );
  OAI22X1TF U155 ( .A0(N686), .A1(N189), .B0(N654), .B1(N186), .Y(N1040) );
  AND2X2TF U156 ( .A(N1012), .B(N1022), .Y(N1013) );
  CLKBUFX2TF U157 ( .A(N584), .Y(N171) );
  OR2X2TF U158 ( .A(N1017), .B(N537), .Y(N844) );
  AND2X2TF U159 ( .A(N1012), .B(N1680), .Y(N188) );
  AND2X2TF U160 ( .A(N1018), .B(N1680), .Y(N182) );
  AND2X2TF U161 ( .A(N1023), .B(N1680), .Y(N185) );
  AND2X2TF U162 ( .A(\OPER1_R1[2] ), .B(N169), .Y(N179) );
  AND2X2TF U163 ( .A(OPER3_R3[2]), .B(N887), .Y(N1185) );
  AND2X2TF U164 ( .A(N243), .B(N278), .Y(N1174) );
  AND2X2TF U165 ( .A(N243), .B(N255), .Y(N1172) );
  AOI32X1TF U166 ( .A0(N555), .A1(N556), .A2(N417), .B0(N553), .B1(N556), .Y(
        N584) );
  CLKINVX1TF U167 ( .A(N335), .Y(N328) );
  ADDFHX2TF U168 ( .A(N423), .B(REG_A[4]), .CI(SUB_X_285_4_N13), .CO(
        SUB_X_285_4_N12), .S(N508) );
  NOR2X4TF U169 ( .A(N1006), .B(N882), .Y(N407) );
  NAND3BXLTF U170 ( .AN(N884), .B(N1005), .C(N1006), .Y(N288) );
  NAND2X1TF U171 ( .A(CODE_TYPE[2]), .B(N555), .Y(N882) );
  ADDFHX2TF U172 ( .A(N230), .B(REG_A[3]), .CI(SUB_X_285_4_N14), .CO(
        SUB_X_285_4_N13), .S(N507) );
  OAI32X1TF U173 ( .A0(STATE[1]), .A1(STATE[3]), .A2(N554), .B0(N733), .B1(
        N207), .Y(N110) );
  CLKINVX2TF U174 ( .A(N399), .Y(N173) );
  OR2X1TF U175 ( .A(N43), .B(N770), .Y(N229) );
  INVX2TF U176 ( .A(N1187), .Y(N172) );
  AND2X2TF U177 ( .A(N193), .B(N1129), .Y(N826) );
  NAND2XLTF U178 ( .A(STATE[1]), .B(N203), .Y(N536) );
  NAND4XLTF U179 ( .A(N554), .B(N671), .C(N670), .D(N669), .Y(N725) );
  NAND2XLTF U180 ( .A(STATE[0]), .B(N207), .Y(N722) );
  INVX2TF U181 ( .A(N141), .Y(N142) );
  INVX2TF U182 ( .A(N869), .Y(N143) );
  INVX2TF U183 ( .A(N826), .Y(N144) );
  INVX2TF U184 ( .A(N826), .Y(N145) );
  INVX2TF U185 ( .A(N1174), .Y(N146) );
  INVX2TF U186 ( .A(N1174), .Y(N147) );
  INVX2TF U187 ( .A(N1172), .Y(N148) );
  INVX2TF U188 ( .A(N1172), .Y(N149) );
  INVX2TF U189 ( .A(N44), .Y(N150) );
  INVX2TF U190 ( .A(N44), .Y(N151) );
  INVX2TF U191 ( .A(N1049), .Y(N152) );
  INVX2TF U192 ( .A(N1049), .Y(N153) );
  INVX2TF U193 ( .A(N1164), .Y(N154) );
  INVX2TF U194 ( .A(N1164), .Y(N155) );
  INVX2TF U195 ( .A(N844), .Y(N156) );
  INVX2TF U196 ( .A(N844), .Y(N157) );
  INVX2TF U197 ( .A(N1165), .Y(N159) );
  INVX2TF U198 ( .A(N1165), .Y(N160) );
  INVX2TF U199 ( .A(N1166), .Y(N161) );
  INVX2TF U200 ( .A(N1166), .Y(N162) );
  INVX2TF U201 ( .A(N163), .Y(N164) );
  INVX2TF U202 ( .A(N163), .Y(N165) );
  INVX2TF U203 ( .A(N1185), .Y(N1660) );
  INVX2TF U204 ( .A(N1185), .Y(N1670) );
  INVX2TF U205 ( .A(N1159), .Y(N1680) );
  INVX2TF U206 ( .A(N1159), .Y(N169) );
  INVX2TF U207 ( .A(N1159), .Y(N170) );
  AOI22XLTF U208 ( .A0(N332), .A1(N849), .B0(N749), .B1(N847), .Y(N291) );
  NOR3X2TF U209 ( .A(N736), .B(N236), .C(\OPER1_R1[2] ), .Y(N1012) );
  AOI22X2TF U210 ( .A0(REG_C[11]), .A1(N583), .B0(N585), .B1(D_DATAIN[3]), .Y(
        N697) );
  AOI22X2TF U211 ( .A0(REG_C[12]), .A1(N583), .B0(N585), .B1(D_DATAIN[4]), .Y(
        N698) );
  AOI22X2TF U212 ( .A0(REG_C[10]), .A1(N583), .B0(N585), .B1(D_DATAIN[2]), .Y(
        N696) );
  AOI22X2TF U213 ( .A0(REG_C[9]), .A1(N583), .B0(N585), .B1(D_DATAIN[1]), .Y(
        N695) );
  AOI22X2TF U214 ( .A0(D_ADDR[5]), .A1(N559), .B0(N558), .B1(D_DATAIN[4]), .Y(
        N577) );
  AOI22X2TF U215 ( .A0(D_ADDR[1]), .A1(N559), .B0(N558), .B1(D_DATAIN[0]), .Y(
        N573) );
  AOI22X2TF U216 ( .A0(D_ADDR[2]), .A1(N559), .B0(N558), .B1(D_DATAIN[1]), .Y(
        N574) );
  AOI22X2TF U217 ( .A0(D_ADDR[4]), .A1(N559), .B0(N558), .B1(D_DATAIN[3]), .Y(
        N576) );
  AOI32X1TF U218 ( .A0(N223), .A1(N231), .A2(N728), .B0(STATE[0]), .B1(N536), 
        .Y(N166) );
  NOR2BX2TF U219 ( .AN(CODE_TYPE[4]), .B(CODE_TYPE[3]), .Y(N417) );
  OAI22X2TF U220 ( .A0(N545), .A1(N557), .B0(N733), .B1(N728), .Y(N715) );
  NOR3X4TF U221 ( .A(N572), .B(N571), .C(N566), .Y(N568) );
  NOR3X4TF U222 ( .A(N572), .B(N571), .C(N594), .Y(N693) );
  NOR3X4TF U223 ( .A(N571), .B(N236), .C(N594), .Y(N593) );
  OAI22XLTF U224 ( .A0(N636), .A1(N191), .B0(N668), .B1(N1177), .Y(N907) );
  OAI211XLTF U225 ( .A0(N735), .A1(N723), .B0(N722), .C0(N1190), .Y(
        NEXT_STATE[0]) );
  NOR3X4TF U226 ( .A(N223), .B(N231), .C(N735), .Y(N558) );
  NAND2X2TF U227 ( .A(N554), .B(STATE[1]), .Y(N735) );
  OAI22XLTF U228 ( .A0(N620), .A1(N1660), .B0(N652), .B1(N1180), .Y(N906) );
  OAI22XLTF U229 ( .A0(N615), .A1(N1660), .B0(N647), .B1(N1180), .Y(N902) );
  OAI22XLTF U230 ( .A0(N613), .A1(N1660), .B0(N645), .B1(N1180), .Y(N890) );
  INVX2TF U231 ( .A(N1190), .Y(N174) );
  INVX2TF U232 ( .A(N845), .Y(N175) );
  NOR2X1TF U233 ( .A(N1006), .B(N1032), .Y(N410) );
  CLKBUFX2TF U234 ( .A(N1170), .Y(N176) );
  CLKBUFX2TF U235 ( .A(N1162), .Y(N177) );
  NOR2BX2TF U236 ( .AN(N1680), .B(N1020), .Y(N1162) );
  CLKBUFX2TF U237 ( .A(N1175), .Y(N178) );
  OAI31X4TF U238 ( .A0(N1017), .A1(N1016), .A2(N1015), .B0(N1014), .Y(N1049)
         );
  NOR2X4TF U239 ( .A(N193), .B(N1129), .Y(N746) );
  NOR3X4TF U240 ( .A(N861), .B(REG_B[3]), .C(N43), .Y(N854) );
  INVX2TF U241 ( .A(N179), .Y(N180) );
  INVX2TF U242 ( .A(N179), .Y(N181) );
  INVX2TF U243 ( .A(N182), .Y(N183) );
  INVX2TF U244 ( .A(N182), .Y(N184) );
  INVX2TF U245 ( .A(N185), .Y(N186) );
  INVX2TF U246 ( .A(N185), .Y(N187) );
  OAI21X2TF U247 ( .A0(N883), .A1(N910), .B0(N1014), .Y(N1128) );
  OAI211X1TF U248 ( .A0(CODE_TYPE[3]), .A1(N876), .B0(N1014), .C0(N206), .Y(
        N885) );
  INVX2TF U249 ( .A(N188), .Y(N189) );
  INVX2TF U250 ( .A(N188), .Y(N190) );
  CLKBUFX2TF U251 ( .A(N1178), .Y(N191) );
  OAI22XLTF U252 ( .A0(N635), .A1(N1178), .B0(N667), .B1(N1177), .Y(N899) );
  OAI22XLTF U253 ( .A0(N640), .A1(N1178), .B0(N672), .B1(N1177), .Y(N912) );
  NOR3X4TF U254 ( .A(N571), .B(N236), .C(N566), .Y(N565) );
  CLKBUFX2TF U255 ( .A(N1173), .Y(N192) );
  NOR2X1TF U256 ( .A(N250), .B(N1118), .Y(N1173) );
  AOI2BB2X2TF U257 ( .B0(D_DATAIN[5]), .B1(N585), .A0N(N421), .A1N(N171), .Y(
        N699) );
  AOI2BB2X2TF U258 ( .B0(D_DATAIN[7]), .B1(N585), .A0N(N414), .A1N(N171), .Y(
        N612) );
  AOI2BB2X2TF U259 ( .B0(D_DATAIN[6]), .B1(N585), .A0N(N416), .A1N(N171), .Y(
        N701) );
  AOI22X2TF U260 ( .A0(REG_C[8]), .A1(N583), .B0(N585), .B1(D_DATAIN[0]), .Y(
        N694) );
  NOR3X4TF U261 ( .A(N210), .B(N877), .C(N878), .Y(N585) );
  AOI22X2TF U262 ( .A0(D_ADDR[7]), .A1(N559), .B0(N558), .B1(D_DATAIN[6]), .Y(
        N579) );
  AOI22X2TF U263 ( .A0(D_ADDR[6]), .A1(N559), .B0(N558), .B1(D_DATAIN[5]), .Y(
        N578) );
  AOI22X2TF U264 ( .A0(D_ADDR[8]), .A1(N559), .B0(N558), .B1(D_DATAIN[7]), .Y(
        N581) );
  AOI22X2TF U265 ( .A0(D_ADDR[3]), .A1(N559), .B0(N558), .B1(D_DATAIN[2]), .Y(
        N575) );
  NOR3X4TF U266 ( .A(N223), .B(N735), .C(STATE[0]), .Y(N559) );
  XOR2X1TF U267 ( .A(REG_A[0]), .B(REG_B[0]), .Y(N504) );
  NAND2BX1TF U268 ( .AN(REG_A[0]), .B(REG_B[0]), .Y(SUB_X_285_4_N16) );
  CMPR32X2TF U269 ( .A(N408), .B(REG_A[10]), .C(SUB_X_285_4_N7), .CO(
        SUB_X_285_4_N6), .S(N514) );
  CMPR32X2TF U270 ( .A(N418), .B(REG_A[9]), .C(SUB_X_285_4_N8), .CO(
        SUB_X_285_4_N7), .S(N513) );
  ADDFHX2TF U271 ( .A(N140), .B(REG_A[2]), .CI(SUB_X_285_4_N15), .CO(
        SUB_X_285_4_N14), .S(N506) );
  XOR2X2TF U272 ( .A(N376), .B(N375), .Y(N381) );
  AOI21X4TF U273 ( .A0(N482), .A1(N245), .B0(N284), .Y(N396) );
  OAI2BB1X4TF U274 ( .A0N(N348), .A1N(N485), .B0(N301), .Y(N376) );
  CLKINVX4TF U275 ( .A(N376), .Y(N373) );
  AOI211X2TF U276 ( .A0(N519), .A1(N244), .B0(N300), .C0(N299), .Y(N301) );
  OA22X1TF U277 ( .A0(N392), .A1(N147), .B0(N393), .B1(N148), .Y(N1119) );
  CLKXOR2X2TF U278 ( .A(N397), .B(N374), .Y(N375) );
  AO21X1TF U279 ( .A0(N341), .A1(N422), .B0(N143), .Y(N5090) );
  NOR2X2TF U280 ( .A(N205), .B(N210), .Y(N1034) );
  AO21X1TF U281 ( .A0(IO_DATAINA[9]), .A1(N192), .B0(N371), .Y(N4720) );
  CLKBUFX2TF U282 ( .A(N348), .Y(N245) );
  CLKBUFX2TF U283 ( .A(N44), .Y(N247) );
  INVX2TF U284 ( .A(N139), .Y(N251) );
  NAND2X1TF U285 ( .A(N205), .B(N250), .Y(N878) );
  NAND2X1TF U286 ( .A(N225), .B(N570), .Y(N566) );
  OAI2BB1X1TF U287 ( .A0N(N245), .A1N(N478), .B0(N347), .Y(N368) );
  NOR3X1TF U288 ( .A(N569), .B(N250), .C(N205), .Y(N876) );
  CLKBUFX2TF U289 ( .A(N399), .Y(N243) );
  AOI211XLTF U290 ( .A0(STATE[0]), .A1(N730), .B0(N243), .C0(N729), .Y(N731)
         );
  AOI31X1TF U291 ( .A0(N42), .A1(N419), .A2(N1004), .B0(N557), .Y(N727) );
  NAND2X1TF U292 ( .A(N5880), .B(N225), .Y(N594) );
  OAI2BB2X1TF U293 ( .B0(N557), .B1(N171), .A0N(N585), .A1N(N558), .Y(N570) );
  AOI21X2TF U294 ( .A0(N484), .A1(N348), .B0(N287), .Y(N395) );
  CLKBUFX2TF U295 ( .A(N865), .Y(N244) );
  OR2X2TF U296 ( .A(N267), .B(N266), .Y(N348) );
  NAND2X1TF U297 ( .A(N1014), .B(N1015), .Y(N1025) );
  NOR2X1TF U298 ( .A(N885), .B(N910), .Y(N887) );
  NOR2X1TF U299 ( .A(N736), .B(N572), .Y(N1018) );
  AOI21X1TF U300 ( .A0(N556), .A1(N171), .B0(N557), .Y(N5880) );
  INVX2TF U301 ( .A(N399), .Y(N1171) );
  INVX2TF U302 ( .A(N863), .Y(N4810) );
  NOR2X2TF U303 ( .A(CODE_TYPE[3]), .B(CODE_TYPE[4]), .Y(N1004) );
  NAND2X1TF U304 ( .A(N205), .B(N210), .Y(N1011) );
  NOR2X2TF U305 ( .A(N158), .B(N569), .Y(N555) );
  OAI211XLTF U306 ( .A0(IO_CONTROL[4]), .A1(N725), .B0(N724), .C0(STATE[1]), 
        .Y(N732) );
  AOI22XLTF U307 ( .A0(REG_A[5]), .A1(N1049), .B0(IO_CONTROL[5]), .B1(N1164), 
        .Y(N1028) );
  NAND2X1TF U308 ( .A(N1014), .B(N1016), .Y(N1024) );
  NAND2X1TF U309 ( .A(N288), .B(N243), .Y(N1186) );
  NAND3X2TF U310 ( .A(N885), .B(N1128), .C(N1151), .Y(N1179) );
  INVX2TF U311 ( .A(N875), .Y(N1014) );
  INVX2TF U312 ( .A(N1190), .Y(N1192) );
  NAND3X1TF U313 ( .A(N203), .B(N207), .C(N724), .Y(N1190) );
  INVX2TF U314 ( .A(N1187), .Y(N1188) );
  NOR2X2TF U315 ( .A(N5890), .B(N594), .Y(N591) );
  NOR2X2TF U316 ( .A(N5890), .B(N566), .Y(N563) );
  INVX2TF U317 ( .A(N559), .Y(N557) );
  OAI211X1TF U318 ( .A0(STATE[1]), .A1(N733), .B0(I_ADDR[0]), .C0(N875), .Y(
        N550) );
  INVX2TF U319 ( .A(N1004), .Y(N877) );
  NAND2X2TF U320 ( .A(N866), .B(N851), .Y(N833) );
  NAND3X1TF U321 ( .A(N417), .B(N1034), .C(N243), .Y(N1118) );
  NAND3X2TF U322 ( .A(N250), .B(N1034), .C(N1004), .Y(N861) );
  NAND2X1TF U323 ( .A(N1004), .B(N876), .Y(N427) );
  NOR2X1TF U324 ( .A(N219), .B(N206), .Y(N1008) );
  OR3X1TF U325 ( .A(N555), .B(N205), .C(CODE_TYPE[3]), .Y(N552) );
  AND2X2TF U326 ( .A(N554), .B(N253), .Y(N399) );
  NOR3BX1TF U327 ( .AN(STATE[0]), .B(STATE[3]), .C(STATE[1]), .Y(N253) );
  OAI32XLTF U328 ( .A0(N231), .A1(STATE[1]), .A2(N554), .B0(N735), .B1(N231), 
        .Y(NEXT_STATE[3]) );
  NOR2XLTF U329 ( .A(STATE[1]), .B(N203), .Y(N734) );
  AO22X1TF U330 ( .A0(N394), .A1(CF_BUF), .B0(N1186), .B1(CF), .Y(N5180) );
  AOI22XLTF U331 ( .A0(REG_A[6]), .A1(N1049), .B0(IO_CONTROL[6]), .B1(N1164), 
        .Y(N1039) );
  NOR2BX1TF U332 ( .AN(N402), .B(N1024), .Y(N1019) );
  NAND2X1TF U333 ( .A(N717), .B(I_ADDR[8]), .Y(N726) );
  NOR2X1TF U334 ( .A(N718), .B(N238), .Y(N717) );
  OAI2BB2XLTF U335 ( .B0(N1192), .B1(N42), .A0N(N1192), .A1N(I_DATAIN[4]), .Y(
        N531) );
  OAI2BB2XLTF U336 ( .B0(N1188), .B1(N403), .A0N(N1188), .A1N(I_DATAIN[6]), 
        .Y(N521) );
  OAI2BB2XLTF U337 ( .B0(N1192), .B1(N572), .A0N(N1192), .A1N(I_DATAIN[0]), 
        .Y(N535) );
  OAI2BB2XLTF U338 ( .B0(N1188), .B1(N209), .A0N(N1188), .A1N(I_DATAIN[1]), 
        .Y(N526) );
  OAI2BB2XLTF U339 ( .B0(N1192), .B1(N225), .A0N(N1192), .A1N(I_DATAIN[2]), 
        .Y(N533) );
  OAI2BB2XLTF U340 ( .B0(N1188), .B1(N402), .A0N(N1188), .A1N(I_DATAIN[5]), 
        .Y(N522) );
  OAI2BB2XLTF U341 ( .B0(N1188), .B1(N204), .A0N(N1188), .A1N(I_DATAIN[2]), 
        .Y(N525) );
  OAI2BB2XLTF U342 ( .B0(N1192), .B1(N219), .A0N(N1192), .A1N(I_DATAIN[6]), 
        .Y(N529) );
  OAI2BB2XLTF U343 ( .B0(N1192), .B1(N571), .A0N(N174), .A1N(I_DATAIN[1]), .Y(
        N534) );
  OAI2BB2XLTF U344 ( .B0(N1192), .B1(N205), .A0N(N174), .A1N(I_DATAIN[5]), .Y(
        N530) );
  OAI2BB2XLTF U345 ( .B0(N1188), .B1(N226), .A0N(N172), .A1N(I_DATAIN[0]), .Y(
        N527) );
  NAND4X1TF U346 ( .A(N223), .B(N203), .C(N207), .D(STATE[0]), .Y(N1187) );
  INVX2TF U347 ( .A(N591), .Y(N590) );
  INVX2TF U348 ( .A(N593), .Y(N592) );
  INVX2TF U349 ( .A(N568), .Y(N567) );
  INVX2TF U350 ( .A(N693), .Y(N611) );
  INVX2TF U351 ( .A(N700), .Y(N702) );
  NAND2X2TF U352 ( .A(N570), .B(N1012), .Y(N560) );
  INVX2TF U353 ( .A(N565), .Y(N564) );
  INVX2TF U354 ( .A(N580), .Y(N582) );
  OAI221XLTF U355 ( .A0(N730), .A1(N550), .B0(N735), .B1(N733), .C0(N549), .Y(
        N1002) );
  NAND4X1TF U356 ( .A(N203), .B(N207), .C(STATE[0]), .D(STATE[3]), .Y(N875) );
  NOR2X1TF U357 ( .A(STATE[3]), .B(STATE[0]), .Y(N724) );
  NOR4XLTF U358 ( .A(N741), .B(N723), .C(N203), .D(N877), .Y(N616) );
  OAI221XLTF U359 ( .A0(REG_A[2]), .A1(N139), .B0(N216), .B1(N845), .C0(N157), 
        .Y(N787) );
  OAI221XLTF U360 ( .A0(REG_A[1]), .A1(N139), .B0(N200), .B1(N845), .C0(N157), 
        .Y(N778) );
  INVX2TF U361 ( .A(N410), .Y(N845) );
  NAND2X1TF U362 ( .A(N151), .B(REG_A[10]), .Y(N816) );
  NAND2X1TF U363 ( .A(N151), .B(REG_A[11]), .Y(N766) );
  NAND2X1TF U364 ( .A(N151), .B(REG_A[7]), .Y(N762) );
  NAND2X1TF U365 ( .A(N151), .B(REG_A[8]), .Y(N745) );
  NAND2BX1TF U366 ( .AN(N1006), .B(N257), .Y(N538) );
  NAND2X1TF U367 ( .A(N205), .B(N158), .Y(N1007) );
  NOR3X1TF U368 ( .A(N252), .B(N537), .C(N865), .Y(N539) );
  OAI21X1TF U369 ( .A0(N734), .A1(N733), .B0(N1187), .Y(NEXT_STATE[2]) );
  INVX2TF U370 ( .A(N1186), .Y(N394) );
  OAI21X1TF U371 ( .A0(N623), .A1(N180), .B0(N1031), .Y(N445) );
  AOI211X1TF U372 ( .A0(N1162), .A1(IO_DATAOUTB[5]), .B0(N1030), .C0(N1029), 
        .Y(N1031) );
  OAI21X1TF U373 ( .A0(N626), .A1(N180), .B0(N1065), .Y(N462) );
  AOI211X1TF U374 ( .A0(N1162), .A1(IO_DATAOUTB[2]), .B0(N1064), .C0(N1063), 
        .Y(N1065) );
  OAI21X1TF U375 ( .A0(N624), .A1(N180), .B0(N1048), .Y(N453) );
  AOI211X1TF U376 ( .A0(N1162), .A1(IO_DATAOUTB[4]), .B0(N1047), .C0(N1046), 
        .Y(N1048) );
  OAI21X1TF U377 ( .A0(N620), .A1(N180), .B0(N1055), .Y(N457) );
  AOI211X1TF U378 ( .A0(N1162), .A1(IO_DATAOUTB[8]), .B0(N1054), .C0(N1053), 
        .Y(N1055) );
  OAI21X1TF U379 ( .A0(N619), .A1(N180), .B0(N1079), .Y(N4700) );
  AOI211X1TF U380 ( .A0(N1162), .A1(IO_DATAOUTB[9]), .B0(N1078), .C0(N1077), 
        .Y(N1079) );
  OAI21X1TF U381 ( .A0(N622), .A1(N180), .B0(N1042), .Y(N449) );
  AOI211X1TF U382 ( .A0(N1162), .A1(IO_DATAOUTB[6]), .B0(N1041), .C0(N1040), 
        .Y(N1042) );
  OAI21X1TF U383 ( .A0(N627), .A1(N180), .B0(N1117), .Y(N489) );
  AOI211X1TF U384 ( .A0(N1162), .A1(IO_DATAOUTB[1]), .B0(N1116), .C0(N1115), 
        .Y(N1117) );
  OAI22X1TF U385 ( .A0(N170), .A1(N609), .B0(N675), .B1(N184), .Y(N1116) );
  OAI21X1TF U386 ( .A0(N613), .A1(N180), .B0(N1127), .Y(N493) );
  AOI211X1TF U387 ( .A0(N177), .A1(N242), .B0(N1126), .C0(N1125), .Y(N1127) );
  OAI22X1TF U388 ( .A0(N169), .A1(N595), .B0(N661), .B1(N184), .Y(N1126) );
  OAI21X1TF U389 ( .A0(N625), .A1(N181), .B0(N1099), .Y(N4800) );
  AOI211X1TF U390 ( .A0(N177), .A1(IO_DATAOUTB[3]), .B0(N1098), .C0(N1097), 
        .Y(N1099) );
  OAI22X1TF U391 ( .A0(N170), .A1(N607), .B0(N673), .B1(N184), .Y(N1098) );
  OAI21X1TF U392 ( .A0(N6160), .A1(N181), .B0(N1150), .Y(N503) );
  AOI211X1TF U393 ( .A0(N177), .A1(IO_DATAOUTB[12]), .B0(N1149), .C0(N1148), 
        .Y(N1150) );
  OAI22X1TF U394 ( .A0(N169), .A1(N598), .B0(N664), .B1(N184), .Y(N1149) );
  OAI21X1TF U395 ( .A0(N618), .A1(N181), .B0(N1089), .Y(N4750) );
  AOI211X1TF U396 ( .A0(N177), .A1(IO_DATAOUTB[10]), .B0(N1088), .C0(N1087), 
        .Y(N1089) );
  OAI22X1TF U397 ( .A0(N170), .A1(N600), .B0(N666), .B1(N184), .Y(N1088) );
  OAI21X1TF U398 ( .A0(N621), .A1(N181), .B0(N739), .Y(N433) );
  AOI211X1TF U399 ( .A0(N177), .A1(IO_DATAOUTB[7]), .B0(N738), .C0(N737), .Y(
        N739) );
  OAI22X1TF U400 ( .A0(N169), .A1(N603), .B0(N669), .B1(N184), .Y(N738) );
  OAI21X1TF U401 ( .A0(N628), .A1(N181), .B0(N1139), .Y(N498) );
  AOI211X1TF U402 ( .A0(N177), .A1(IO_DATAOUTB[0]), .B0(N1138), .C0(N1137), 
        .Y(N1139) );
  OAI22X1TF U403 ( .A0(N170), .A1(N610), .B0(N676), .B1(N184), .Y(N1138) );
  OAI21X1TF U404 ( .A0(N614), .A1(N181), .B0(N1107), .Y(N4840) );
  AOI211X1TF U405 ( .A0(N177), .A1(N241), .B0(N1106), .C0(N1105), .Y(N1107) );
  OAI22X1TF U406 ( .A0(N169), .A1(N596), .B0(N662), .B1(N184), .Y(N1106) );
  OAI21X1TF U407 ( .A0(N615), .A1(N181), .B0(N1073), .Y(N466) );
  AOI211X1TF U408 ( .A0(N177), .A1(N240), .B0(N1072), .C0(N1071), .Y(N1073) );
  OAI22X1TF U409 ( .A0(N170), .A1(N597), .B0(N663), .B1(N184), .Y(N1072) );
  OAI21X1TF U410 ( .A0(N617), .A1(N181), .B0(N1163), .Y(N5080) );
  AOI211X1TF U411 ( .A0(N177), .A1(IO_DATAOUTB[11]), .B0(N1161), .C0(N1160), 
        .Y(N1163) );
  OAI22X1TF U412 ( .A0(N169), .A1(N599), .B0(N665), .B1(N184), .Y(N1161) );
  OAI21X1TF U413 ( .A0(N1170), .A1(N691), .B0(N1114), .Y(N488) );
  AOI211X1TF U414 ( .A0(IO_DATAOUTB[1]), .A1(N164), .B0(N1113), .C0(N1112), 
        .Y(N1114) );
  OAI21X1TF U415 ( .A0(N1170), .A1(N678), .B0(N1104), .Y(N4830) );
  AOI211X1TF U416 ( .A0(N241), .A1(N164), .B0(N1103), .C0(N1102), .Y(N1104) );
  OAI21X1TF U417 ( .A0(N1170), .A1(N681), .B0(N1158), .Y(N5070) );
  AOI211X1TF U418 ( .A0(IO_DATAOUTB[11]), .A1(N165), .B0(N1157), .C0(N1156), 
        .Y(N1158) );
  OAI21X1TF U419 ( .A0(N1170), .A1(N677), .B0(N1124), .Y(N492) );
  AOI211X1TF U420 ( .A0(N242), .A1(N165), .B0(N1123), .C0(N1122), .Y(N1124) );
  OAI21X1TF U421 ( .A0(N1170), .A1(N680), .B0(N1147), .Y(N502) );
  AOI211X1TF U422 ( .A0(IO_DATAOUTB[12]), .A1(N165), .B0(N1146), .C0(N1145), 
        .Y(N1147) );
  OAI21X1TF U423 ( .A0(N1170), .A1(N679), .B0(N1070), .Y(N465) );
  AOI211X1TF U424 ( .A0(N240), .A1(N165), .B0(N1069), .C0(N1068), .Y(N1070) );
  OAI21X1TF U425 ( .A0(N176), .A1(N690), .B0(N1062), .Y(N461) );
  AOI211X1TF U426 ( .A0(IO_DATAOUTB[2]), .A1(N164), .B0(N1061), .C0(N1060), 
        .Y(N1062) );
  OAI21X1TF U427 ( .A0(N176), .A1(N685), .B0(N1169), .Y(N5110) );
  AOI211X1TF U428 ( .A0(IO_DATAOUTB[7]), .A1(N164), .B0(N1168), .C0(N1167), 
        .Y(N1169) );
  OAI21X1TF U429 ( .A0(N176), .A1(N682), .B0(N1086), .Y(N4740) );
  AOI211X1TF U430 ( .A0(IO_DATAOUTB[10]), .A1(N164), .B0(N1085), .C0(N1084), 
        .Y(N1086) );
  OAI21X1TF U431 ( .A0(N176), .A1(N683), .B0(N1076), .Y(N469) );
  AOI211X1TF U432 ( .A0(IO_DATAOUTB[9]), .A1(N164), .B0(N1075), .C0(N1074), 
        .Y(N1076) );
  OAI21X1TF U433 ( .A0(N176), .A1(N689), .B0(N1096), .Y(N4790) );
  AOI211X1TF U434 ( .A0(IO_DATAOUTB[3]), .A1(N164), .B0(N1095), .C0(N1094), 
        .Y(N1096) );
  OAI21X1TF U435 ( .A0(N176), .A1(N684), .B0(N1052), .Y(N456) );
  AOI211X1TF U436 ( .A0(IO_DATAOUTB[8]), .A1(N164), .B0(N1051), .C0(N1050), 
        .Y(N1052) );
  OAI21X1TF U437 ( .A0(N176), .A1(N692), .B0(N1136), .Y(N497) );
  AOI211X1TF U438 ( .A0(IO_DATAOUTB[0]), .A1(N165), .B0(N1135), .C0(N1134), 
        .Y(N1136) );
  OAI21X1TF U439 ( .A0(N420), .A1(N53), .B0(N909), .Y(N440) );
  NOR3X1TF U440 ( .A(N908), .B(N907), .C(N906), .Y(N909) );
  OAI22X1TF U441 ( .A0(N684), .A1(N1175), .B0(N226), .B1(N1151), .Y(N908) );
  OAI21X1TF U442 ( .A0(N415), .A1(N1179), .B0(N897), .Y(N437) );
  NOR3X1TF U443 ( .A(N896), .B(N895), .C(N894), .Y(N897) );
  OAI22X1TF U444 ( .A0(N678), .A1(N1175), .B0(N403), .B1(N1151), .Y(N896) );
  OAI21X1TF U445 ( .A0(N413), .A1(N53), .B0(N905), .Y(N439) );
  NOR3X1TF U446 ( .A(N904), .B(N903), .C(N902), .Y(N905) );
  OAI22X1TF U447 ( .A0(N679), .A1(N1175), .B0(N402), .B1(N1151), .Y(N904) );
  OAI21X1TF U448 ( .A0(N412), .A1(N53), .B0(N893), .Y(N436) );
  NOR3X1TF U449 ( .A(N892), .B(N891), .C(N890), .Y(N893) );
  OAI22X1TF U450 ( .A0(N677), .A1(N1175), .B0(N404), .B1(N1151), .Y(N892) );
  OAI211X1TF U451 ( .A0(N1170), .A1(N687), .B0(N1028), .C0(N1027), .Y(N444) );
  AOI21X1TF U452 ( .A0(IO_DATAOUTB[5]), .A1(N165), .B0(N1026), .Y(N1027) );
  OAI211X1TF U453 ( .A0(N1170), .A1(N686), .B0(N1039), .C0(N1038), .Y(N448) );
  AOI21X1TF U454 ( .A0(IO_DATAOUTB[6]), .A1(N165), .B0(N1037), .Y(N1038) );
  OAI211X1TF U455 ( .A0(N1170), .A1(N688), .B0(N1045), .C0(N1044), .Y(N452) );
  AOI21X1TF U456 ( .A0(IO_DATAOUTB[4]), .A1(N165), .B0(N1043), .Y(N1044) );
  NOR2X1TF U457 ( .A(N571), .B(N236), .Y(N1023) );
  NOR2X1TF U458 ( .A(N1024), .B(N402), .Y(N1021) );
  AOI22X1TF U459 ( .A0(REG_A[4]), .A1(N1049), .B0(IO_CONTROL[4]), .B1(N1164), 
        .Y(N1045) );
  AOI31X4TF U460 ( .A0(N403), .A1(N401), .A2(N1019), .B0(N1013), .Y(N1170) );
  INVX2TF U461 ( .A(N1025), .Y(N1022) );
  OAI211X1TF U462 ( .A0(N219), .A1(N1011), .B0(N1010), .C0(N1009), .Y(N1015)
         );
  AOI32X1TF U463 ( .A0(N417), .A1(N257), .A2(N569), .B0(N1008), .B1(N1007), 
        .Y(N1010) );
  OAI21X1TF U464 ( .A0(N628), .A1(N1670), .B0(N1133), .Y(N496) );
  NOR3X1TF U465 ( .A(N1132), .B(N1131), .C(N1130), .Y(N1133) );
  OAI22X1TF U466 ( .A0(N660), .A1(N249), .B0(N1129), .B1(N1179), .Y(N1130) );
  OAI22X1TF U467 ( .A0(N644), .A1(N1178), .B0(N676), .B1(N248), .Y(N1131) );
  OAI22X1TF U468 ( .A0(N692), .A1(N1175), .B0(N226), .B1(N1128), .Y(N1132) );
  OAI21X1TF U469 ( .A0(N627), .A1(N1670), .B0(N1111), .Y(N487) );
  NOR3X1TF U470 ( .A(N1110), .B(N1109), .C(N1108), .Y(N1111) );
  OAI22X1TF U471 ( .A0(N659), .A1(N249), .B0(N193), .B1(N1179), .Y(N1108) );
  OAI22X1TF U472 ( .A0(N643), .A1(N1178), .B0(N675), .B1(N248), .Y(N1109) );
  OAI22X1TF U473 ( .A0(N691), .A1(N1175), .B0(N209), .B1(N1128), .Y(N1110) );
  OAI21X1TF U474 ( .A0(N624), .A1(N1670), .B0(N914), .Y(N441) );
  NOR3X1TF U475 ( .A(N913), .B(N912), .C(N911), .Y(N914) );
  OAI22X1TF U476 ( .A0(N656), .A1(N249), .B0(N423), .B1(N1179), .Y(N911) );
  OAI22X1TF U477 ( .A0(N688), .A1(N178), .B0(N401), .B1(N1176), .Y(N913) );
  OAI21X1TF U478 ( .A0(N622), .A1(N1670), .B0(N918), .Y(N442) );
  NOR3X1TF U479 ( .A(N917), .B(N916), .C(N915), .Y(N918) );
  OAI22X1TF U480 ( .A0(N654), .A1(N249), .B0(N406), .B1(N1179), .Y(N915) );
  OAI22X1TF U481 ( .A0(N638), .A1(N1178), .B0(N670), .B1(N248), .Y(N916) );
  OAI22X1TF U482 ( .A0(N686), .A1(N178), .B0(N403), .B1(N1176), .Y(N917) );
  OAI21X1TF U483 ( .A0(N625), .A1(N1670), .B0(N1093), .Y(N4780) );
  NOR3X1TF U484 ( .A(N1092), .B(N1091), .C(N1090), .Y(N1093) );
  OAI22X1TF U485 ( .A0(N657), .A1(N249), .B0(N230), .B1(N1179), .Y(N1090) );
  OAI22X1TF U486 ( .A0(N641), .A1(N1178), .B0(N673), .B1(N248), .Y(N1091) );
  OAI22X1TF U487 ( .A0(N689), .A1(N1175), .B0(N400), .B1(N1128), .Y(N1092) );
  OAI21X1TF U488 ( .A0(N621), .A1(N1670), .B0(N1184), .Y(N5140) );
  NOR3X1TF U489 ( .A(N1183), .B(N1182), .C(N1181), .Y(N1184) );
  OAI22X1TF U490 ( .A0(N653), .A1(N249), .B0(N405), .B1(N1179), .Y(N1181) );
  OAI22X1TF U491 ( .A0(N637), .A1(N1178), .B0(N669), .B1(N248), .Y(N1182) );
  OAI22X1TF U492 ( .A0(N404), .A1(N1176), .B0(N685), .B1(N1175), .Y(N1183) );
  OAI21X1TF U493 ( .A0(N623), .A1(N1670), .B0(N1003), .Y(N443) );
  NOR3X1TF U494 ( .A(N921), .B(N920), .C(N919), .Y(N1003) );
  OAI22X1TF U495 ( .A0(N655), .A1(N249), .B0(N424), .B1(N1179), .Y(N919) );
  OAI22X1TF U496 ( .A0(N639), .A1(N1178), .B0(N671), .B1(N248), .Y(N920) );
  OAI22X1TF U497 ( .A0(N687), .A1(N178), .B0(N402), .B1(N1176), .Y(N921) );
  OAI21X1TF U498 ( .A0(N409), .A1(N53), .B0(N1155), .Y(N5060) );
  NOR3X1TF U499 ( .A(N1154), .B(N1153), .C(N1152), .Y(N1155) );
  OAI22X1TF U500 ( .A0(N617), .A1(N1660), .B0(N649), .B1(N1180), .Y(N1152) );
  OAI22X1TF U501 ( .A0(N633), .A1(N191), .B0(N665), .B1(N248), .Y(N1153) );
  OAI22X1TF U502 ( .A0(N681), .A1(N178), .B0(N400), .B1(N1151), .Y(N1154) );
  OAI21X1TF U503 ( .A0(N411), .A1(N53), .B0(N1144), .Y(N501) );
  NOR3X1TF U504 ( .A(N1143), .B(N1142), .C(N1141), .Y(N1144) );
  OAI22X1TF U505 ( .A0(N6160), .A1(N1670), .B0(N648), .B1(N1180), .Y(N1141) );
  OAI22X1TF U506 ( .A0(N632), .A1(N191), .B0(N664), .B1(N248), .Y(N1142) );
  OAI22X1TF U507 ( .A0(N680), .A1(N178), .B0(N401), .B1(N1151), .Y(N1143) );
  OAI21X1TF U508 ( .A0(N626), .A1(N1670), .B0(N1059), .Y(N460) );
  NOR3X1TF U509 ( .A(N1058), .B(N1057), .C(N1056), .Y(N1059) );
  OAI22X1TF U510 ( .A0(N658), .A1(N249), .B0(N140), .B1(N1179), .Y(N1056) );
  OAI22X1TF U511 ( .A0(N642), .A1(N191), .B0(N674), .B1(N248), .Y(N1057) );
  OAI22X1TF U512 ( .A0(N690), .A1(N1175), .B0(N204), .B1(N1128), .Y(N1058) );
  OAI21X1TF U513 ( .A0(N418), .A1(N53), .B0(N901), .Y(N438) );
  NOR3X1TF U514 ( .A(N900), .B(N899), .C(N898), .Y(N901) );
  OAI22X1TF U515 ( .A0(N619), .A1(N1660), .B0(N651), .B1(N249), .Y(N898) );
  OAI22X1TF U516 ( .A0(N683), .A1(N178), .B0(N209), .B1(N1151), .Y(N900) );
  OAI21X1TF U517 ( .A0(N408), .A1(N53), .B0(N1083), .Y(N4730) );
  NOR3X1TF U518 ( .A(N1082), .B(N1081), .C(N1080), .Y(N1083) );
  OAI22X1TF U519 ( .A0(N618), .A1(N1660), .B0(N650), .B1(N249), .Y(N1080) );
  NOR2X1TF U520 ( .A(OPER3_R3[0]), .B(N888), .Y(N889) );
  OAI22X1TF U521 ( .A0(N634), .A1(N1178), .B0(N666), .B1(N248), .Y(N1081) );
  NOR2X1TF U522 ( .A(OPER3_R3[1]), .B(N888), .Y(N886) );
  NAND3X2TF U523 ( .A(OPER3_R3[0]), .B(OPER3_R3[1]), .C(N887), .Y(N1178) );
  OAI22X1TF U524 ( .A0(N682), .A1(N178), .B0(N204), .B1(N1151), .Y(N1082) );
  NAND2X2TF U525 ( .A(N884), .B(N1014), .Y(N1151) );
  AOI211X1TF U526 ( .A0(N741), .A1(N740), .B0(CODE_TYPE[2]), .C0(N1033), .Y(
        N884) );
  OAI211X1TF U527 ( .A0(N882), .A1(N206), .B0(N881), .C0(N880), .Y(N910) );
  INVX2TF U528 ( .A(N1011), .Y(N419) );
  AOI21X1TF U529 ( .A0(N879), .A1(N878), .B0(N877), .Y(N883) );
  AOI21X1TF U530 ( .A0(D_ADDR[2]), .A1(N721), .B0(N704), .Y(N812) );
  OAI21X1TF U531 ( .A0(N715), .A1(N234), .B0(N703), .Y(N704) );
  OAI211X1TF U532 ( .A0(I_ADDR[1]), .A1(I_ADDR[2]), .B0(N712), .C0(N705), .Y(
        N703) );
  AOI211X1TF U533 ( .A0(N721), .A1(D_ADDR[3]), .B0(N707), .C0(N706), .Y(N811)
         );
  AOI211X1TF U534 ( .A0(N705), .A1(N208), .B0(N708), .C0(N716), .Y(N706) );
  NOR2X1TF U535 ( .A(N208), .B(N715), .Y(N707) );
  AOI21X1TF U536 ( .A0(D_ADDR[1]), .A1(N721), .B0(N547), .Y(N860) );
  AOI22X1TF U537 ( .A0(I_ADDR[1]), .A1(N715), .B0(N716), .B1(N224), .Y(N547)
         );
  AOI211X1TF U538 ( .A0(N721), .A1(D_ADDR[7]), .B0(N720), .C0(N719), .Y(N804)
         );
  AOI211X1TF U539 ( .A0(N718), .A1(N238), .B0(N717), .C0(N716), .Y(N719) );
  NOR2X1TF U540 ( .A(N238), .B(N715), .Y(N720) );
  AOI211X1TF U541 ( .A0(N721), .A1(D_ADDR[5]), .B0(N711), .C0(N710), .Y(N809)
         );
  AOI211X1TF U542 ( .A0(N709), .A1(N235), .B0(N713), .C0(N716), .Y(N710) );
  NOR2X1TF U543 ( .A(N235), .B(N715), .Y(N711) );
  OAI32X1TF U544 ( .A0(N548), .A1(N717), .A2(I_ADDR[8]), .B0(N712), .B1(N548), 
        .Y(N859) );
  INVX2TF U545 ( .A(N716), .Y(N712) );
  INVX2TF U546 ( .A(N715), .Y(N714) );
  NOR2X1TF U547 ( .A(N709), .B(N235), .Y(N713) );
  NOR3X1TF U548 ( .A(N224), .B(N234), .C(N208), .Y(N708) );
  NOR2X2TF U549 ( .A(N557), .B(N546), .Y(N721) );
  AOI32X1TF U550 ( .A0(N544), .A1(N1008), .A2(N237), .B0(N543), .B1(N1008), 
        .Y(N546) );
  OAI22X1TF U551 ( .A0(N740), .A1(N237), .B0(N542), .B1(N541), .Y(N543) );
  OAI22X1TF U552 ( .A0(CF), .A1(N879), .B0(N540), .B1(N205), .Y(N541) );
  AOI21X1TF U553 ( .A0(CF), .A1(N210), .B0(N42), .Y(N540) );
  AOI22X1TF U554 ( .A0(N174), .A1(N1189), .B0(N206), .B1(N1190), .Y(N528) );
  AOI22X1TF U555 ( .A0(N174), .A1(N1191), .B0(N569), .B1(N1190), .Y(N532) );
  AOI22X1TF U556 ( .A0(N172), .A1(N1189), .B0(N404), .B1(N1187), .Y(N520) );
  INVX2TF U557 ( .A(I_DATAIN[7]), .Y(N1189) );
  AOI22X1TF U558 ( .A0(N172), .A1(N1191), .B0(N400), .B1(N1187), .Y(N524) );
  INVX2TF U559 ( .A(I_DATAIN[3]), .Y(N1191) );
  AOI22X1TF U560 ( .A0(N693), .A1(N701), .B0(N630), .B1(N611), .Y(N930) );
  AOI22X1TF U561 ( .A0(N591), .A1(N701), .B0(N662), .B1(N590), .Y(N946) );
  AOI22X1TF U562 ( .A0(N593), .A1(N701), .B0(N646), .B1(N592), .Y(N938) );
  AOI22X1TF U563 ( .A0(N593), .A1(N699), .B0(N647), .B1(N592), .Y(N939) );
  AOI22X1TF U564 ( .A0(N591), .A1(N612), .B0(N661), .B1(N590), .Y(N945) );
  AOI22X1TF U565 ( .A0(N593), .A1(N612), .B0(N645), .B1(N592), .Y(N937) );
  AOI22X1TF U566 ( .A0(N693), .A1(N612), .B0(N629), .B1(N611), .Y(N929) );
  AOI22X1TF U567 ( .A0(N591), .A1(N699), .B0(N663), .B1(N590), .Y(N947) );
  AOI22X1TF U568 ( .A0(N693), .A1(N699), .B0(N631), .B1(N611), .Y(N931) );
  AOI22X1TF U569 ( .A0(N702), .A1(N701), .B0(N614), .B1(N700), .Y(N922) );
  AOI22X1TF U570 ( .A0(N702), .A1(N699), .B0(N615), .B1(N700), .Y(N923) );
  AOI22X1TF U571 ( .A0(N702), .A1(N612), .B0(N613), .B1(N700), .Y(N1001) );
  AOI22X1TF U572 ( .A0(N587), .A1(N699), .B0(N679), .B1(N586), .Y(N955) );
  AOI22X1TF U573 ( .A0(N587), .A1(N612), .B0(N677), .B1(N586), .Y(N953) );
  AOI22X1TF U574 ( .A0(N587), .A1(N701), .B0(N678), .B1(N586), .Y(N954) );
  AOI22X1TF U575 ( .A0(N563), .A1(N581), .B0(N669), .B1(N562), .Y(N985) );
  AOI22X1TF U576 ( .A0(N591), .A1(N694), .B0(N668), .B1(N590), .Y(N952) );
  AOI22X1TF U577 ( .A0(N591), .A1(N697), .B0(N665), .B1(N590), .Y(N949) );
  AOI22X1TF U578 ( .A0(N593), .A1(N694), .B0(N652), .B1(N592), .Y(N944) );
  AOI22X1TF U579 ( .A0(N563), .A1(N575), .B0(N674), .B1(N562), .Y(N990) );
  AOI22X1TF U580 ( .A0(N563), .A1(N579), .B0(N670), .B1(N562), .Y(N986) );
  AOI22X1TF U581 ( .A0(N563), .A1(N578), .B0(N671), .B1(N562), .Y(N987) );
  AOI22X1TF U582 ( .A0(N568), .A1(N579), .B0(N638), .B1(N567), .Y(N970) );
  AOI22X1TF U583 ( .A0(N568), .A1(N578), .B0(N639), .B1(N567), .Y(N971) );
  AOI22X1TF U584 ( .A0(N563), .A1(N577), .B0(N672), .B1(N562), .Y(N988) );
  INVX2TF U585 ( .A(N563), .Y(N562) );
  AOI22X1TF U586 ( .A0(N568), .A1(N581), .B0(N637), .B1(N567), .Y(N969) );
  AOI22X1TF U587 ( .A0(N568), .A1(N575), .B0(N642), .B1(N567), .Y(N974) );
  AOI22X1TF U588 ( .A0(N693), .A1(N694), .B0(N636), .B1(N611), .Y(N936) );
  AOI22X1TF U589 ( .A0(N702), .A1(N698), .B0(N6160), .B1(N700), .Y(N924) );
  AOI22X1TF U590 ( .A0(N702), .A1(N694), .B0(N620), .B1(N700), .Y(N928) );
  AOI22X1TF U591 ( .A0(N702), .A1(N695), .B0(N619), .B1(N700), .Y(N927) );
  AOI22X1TF U592 ( .A0(N702), .A1(N697), .B0(N617), .B1(N700), .Y(N925) );
  AOI22X1TF U593 ( .A0(N702), .A1(N696), .B0(N618), .B1(N700), .Y(N926) );
  NAND4X2TF U594 ( .A(N572), .B(N571), .C(\OPER1_R1[2] ), .D(N5880), .Y(N700)
         );
  AOI22X1TF U595 ( .A0(N587), .A1(N694), .B0(N684), .B1(N586), .Y(N960) );
  AOI22X1TF U596 ( .A0(N587), .A1(N697), .B0(N681), .B1(N586), .Y(N957) );
  AOI22X1TF U597 ( .A0(N587), .A1(N698), .B0(N680), .B1(N586), .Y(N956) );
  AOI22X1TF U598 ( .A0(N587), .A1(N695), .B0(N683), .B1(N586), .Y(N959) );
  AOI22X1TF U599 ( .A0(N587), .A1(N696), .B0(N682), .B1(N586), .Y(N958) );
  INVX2TF U600 ( .A(N171), .Y(N583) );
  INVX2TF U601 ( .A(N586), .Y(N587) );
  NAND2X2TF U602 ( .A(N5880), .B(N1012), .Y(N586) );
  AOI22X1TF U603 ( .A0(N561), .A1(N573), .B0(N692), .B1(N560), .Y(N1000) );
  AOI22X1TF U604 ( .A0(N561), .A1(N578), .B0(N687), .B1(N560), .Y(N995) );
  AOI22X1TF U605 ( .A0(N561), .A1(N576), .B0(N689), .B1(N560), .Y(N997) );
  AOI22X1TF U606 ( .A0(N561), .A1(N575), .B0(N690), .B1(N560), .Y(N998) );
  AOI22X1TF U607 ( .A0(N561), .A1(N579), .B0(N686), .B1(N560), .Y(N994) );
  AOI22X1TF U608 ( .A0(N561), .A1(N574), .B0(N691), .B1(N560), .Y(N999) );
  AOI22X1TF U609 ( .A0(N561), .A1(N577), .B0(N688), .B1(N560), .Y(N996) );
  AOI22X1TF U610 ( .A0(N561), .A1(N581), .B0(N685), .B1(N560), .Y(N993) );
  AOI22X1TF U611 ( .A0(N565), .A1(N581), .B0(N653), .B1(N564), .Y(N977) );
  AOI22X1TF U612 ( .A0(N565), .A1(N579), .B0(N654), .B1(N564), .Y(N978) );
  AOI22X1TF U613 ( .A0(N565), .A1(N576), .B0(N657), .B1(N564), .Y(N981) );
  AOI22X1TF U614 ( .A0(N565), .A1(N578), .B0(N655), .B1(N564), .Y(N979) );
  AOI22X1TF U615 ( .A0(N565), .A1(N575), .B0(N658), .B1(N564), .Y(N982) );
  AOI22X1TF U616 ( .A0(N582), .A1(N579), .B0(N622), .B1(N580), .Y(N962) );
  AOI22X1TF U617 ( .A0(N582), .A1(N578), .B0(N623), .B1(N580), .Y(N963) );
  AOI22X1TF U618 ( .A0(N582), .A1(N581), .B0(N621), .B1(N580), .Y(N961) );
  AOI22X1TF U619 ( .A0(N582), .A1(N575), .B0(N626), .B1(N580), .Y(N966) );
  AOI22X1TF U620 ( .A0(N582), .A1(N576), .B0(N625), .B1(N580), .Y(N965) );
  AOI22X1TF U621 ( .A0(N582), .A1(N573), .B0(N628), .B1(N580), .Y(N968) );
  AOI22X1TF U622 ( .A0(N582), .A1(N577), .B0(N624), .B1(N580), .Y(N964) );
  AOI22X1TF U623 ( .A0(N582), .A1(N574), .B0(N627), .B1(N580), .Y(N967) );
  NAND4X2TF U624 ( .A(N571), .B(N572), .C(\OPER1_R1[2] ), .D(N570), .Y(N580)
         );
  INVX2TF U625 ( .A(N585), .Y(N556) );
  AOI22X1TF U626 ( .A0(I_ADDR[0]), .A1(N595), .B0(N603), .B1(N221), .Y(
        D_DATAOUT[7]) );
  AOI22X1TF U627 ( .A0(I_ADDR[0]), .A1(N596), .B0(N604), .B1(N221), .Y(
        D_DATAOUT[6]) );
  AOI22X1TF U628 ( .A0(I_ADDR[0]), .A1(N597), .B0(N605), .B1(N221), .Y(
        D_DATAOUT[5]) );
  AOI22X1TF U629 ( .A0(I_ADDR[0]), .A1(N598), .B0(N606), .B1(N221), .Y(
        D_DATAOUT[4]) );
  AOI22X1TF U630 ( .A0(I_ADDR[0]), .A1(N599), .B0(N607), .B1(N221), .Y(
        D_DATAOUT[3]) );
  AOI22X1TF U631 ( .A0(I_ADDR[0]), .A1(N600), .B0(N608), .B1(N221), .Y(
        D_DATAOUT[2]) );
  AOI22X1TF U632 ( .A0(I_ADDR[0]), .A1(N601), .B0(N609), .B1(N221), .Y(
        D_DATAOUT[1]) );
  AOI22X1TF U633 ( .A0(I_ADDR[0]), .A1(N602), .B0(N610), .B1(N221), .Y(
        D_DATAOUT[0]) );
  NOR2X1TF U634 ( .A(N243), .B(N558), .Y(N549) );
  INVX2TF U635 ( .A(N724), .Y(N733) );
  AOI21X1TF U636 ( .A0(N363), .A1(N1174), .B0(N362), .Y(N364) );
  AOI22X1TF U637 ( .A0(IO_DATAINB[4]), .A1(N246), .B0(D_ADDR[5]), .B1(N1171), 
        .Y(N360) );
  AOI22X1TF U638 ( .A0(N1140), .A1(IO_STATUS[1]), .B0(N192), .B1(IO_DATAINA[1]), .Y(N1120) );
  AOI22X1TF U639 ( .A0(IO_DATAINB[1]), .A1(N389), .B0(D_ADDR[2]), .B1(N173), 
        .Y(N1121) );
  AOI21X1TF U640 ( .A0(N368), .A1(N1172), .B0(N366), .Y(N367) );
  OAI21X1TF U641 ( .A0(N385), .A1(N146), .B0(N365), .Y(N366) );
  AOI22X1TF U642 ( .A0(IO_DATAINB[8]), .A1(N246), .B0(REG_C[8]), .B1(N1171), 
        .Y(N365) );
  OAI211X1TF U643 ( .A0(N372), .A1(N148), .B0(N370), .C0(N369), .Y(N371) );
  AOI21X1TF U644 ( .A0(N512), .A1(N244), .B0(N346), .Y(N347) );
  OAI21X1TF U645 ( .A0(N831), .A1(N821), .B0(N345), .Y(N346) );
  OAI22X1TF U646 ( .A0(N834), .A1(N835), .B0(N824), .B1(N871), .Y(N343) );
  OAI22X1TF U647 ( .A0(N825), .A1(N833), .B0(N832), .B1(N864), .Y(N823) );
  NOR2X1TF U648 ( .A(N342), .B(N232), .Y(N344) );
  AOI22X1TF U649 ( .A0(REG_A[8]), .A1(N410), .B0(N407), .B1(N232), .Y(N819) );
  AOI22X1TF U650 ( .A0(IO_DATAINB[9]), .A1(N246), .B0(REG_C[9]), .B1(N1171), 
        .Y(N370) );
  AOI21X1TF U651 ( .A0(N479), .A1(N245), .B0(N319), .Y(N372) );
  AOI211X1TF U652 ( .A0(REG_A[9]), .A1(N317), .B0(N813), .C0(N316), .Y(N318)
         );
  OAI21X1TF U653 ( .A0(N806), .A1(N831), .B0(N315), .Y(N316) );
  AOI211X1TF U654 ( .A0(N854), .A1(N839), .B0(N314), .C0(N814), .Y(N315) );
  OAI22X1TF U655 ( .A0(N838), .A1(N833), .B0(N803), .B1(N229), .Y(N814) );
  NOR2X1TF U656 ( .A(N864), .B(N807), .Y(N314) );
  AOI22X1TF U657 ( .A0(REG_A[9]), .A1(N175), .B0(N252), .B1(N212), .Y(N805) );
  AOI21X1TF U658 ( .A0(N481), .A1(N245), .B0(N307), .Y(N383) );
  AOI211X1TF U659 ( .A0(REG_A[11]), .A1(N305), .B0(N304), .C0(N760), .Y(N306)
         );
  AOI22X1TF U660 ( .A0(REG_A[11]), .A1(N410), .B0(N252), .B1(N222), .Y(N757)
         );
  OAI21X1TF U661 ( .A0(N759), .A1(N864), .B0(N303), .Y(N304) );
  AOI211X1TF U662 ( .A0(N758), .A1(N341), .B0(N302), .C0(N761), .Y(N303) );
  OAI22X1TF U663 ( .A0(N794), .A1(N871), .B0(N833), .B1(N797), .Y(N761) );
  NOR2X1TF U664 ( .A(N835), .B(N802), .Y(N302) );
  OAI211X1TF U665 ( .A0(N390), .A1(N149), .B0(N1036), .C0(N1035), .Y(N447) );
  AOI22X1TF U666 ( .A0(IO_DATAINA[5]), .A1(N192), .B0(N1174), .B1(N361), .Y(
        N1035) );
  INVX2TF U667 ( .A(N820), .Y(N824) );
  INVX2TF U668 ( .A(N848), .Y(N825) );
  INVX2TF U669 ( .A(N850), .Y(N834) );
  AOI22X1TF U670 ( .A0(IO_DATAINB[5]), .A1(N389), .B0(D_ADDR[6]), .B1(N173), 
        .Y(N1036) );
  AOI21X1TF U671 ( .A0(N387), .A1(N1174), .B0(N386), .Y(N388) );
  OAI21X1TF U672 ( .A0(N385), .A1(N148), .B0(N384), .Y(N386) );
  AOI22X1TF U673 ( .A0(IO_DATAINB[7]), .A1(N389), .B0(D_ADDR[8]), .B1(N1171), 
        .Y(N384) );
  OAI211X1TF U674 ( .A0(N391), .A1(N147), .B0(N1101), .C0(N11000), .Y(N4820)
         );
  AOI22X1TF U675 ( .A0(IO_DATAINA[3]), .A1(N192), .B0(N1172), .B1(N363), .Y(
        N11000) );
  OAI211X1TF U676 ( .A0(N802), .A1(N837), .B0(N801), .C0(N352), .Y(N363) );
  OAI21X1TF U677 ( .A0(N794), .A1(N831), .B0(N350), .Y(N351) );
  AOI21X1TF U678 ( .A0(N507), .A1(N865), .B0(N349), .Y(N350) );
  AOI211X1TF U679 ( .A0(REG_A[5]), .A1(N151), .B0(N792), .C0(N791), .Y(N793)
         );
  INVX2TF U680 ( .A(N749), .Y(N794) );
  NOR4BX1TF U681 ( .AN(N753), .B(N752), .C(N751), .D(N750), .Y(N795) );
  AOI221X1TF U682 ( .A0(N211), .A1(N407), .B0(REG_A[3]), .B1(N175), .C0(N798), 
        .Y(N799) );
  OAI21X1TF U683 ( .A0(REG_B[3]), .A1(N139), .B0(N796), .Y(N800) );
  AOI211X1TF U684 ( .A0(REG_A[11]), .A1(N422), .B0(N756), .C0(N755), .Y(N802)
         );
  OAI22X1TF U685 ( .A0(N774), .A1(N202), .B0(N247), .B1(N217), .Y(N755) );
  INVX2TF U686 ( .A(N754), .Y(N756) );
  AOI22X1TF U687 ( .A0(IO_DATAINB[3]), .A1(N389), .B0(D_ADDR[4]), .B1(N1171), 
        .Y(N1101) );
  AOI21X1TF U688 ( .A0(N387), .A1(N1172), .B0(N358), .Y(N359) );
  OAI21X1TF U689 ( .A0(N390), .A1(N147), .B0(N357), .Y(N358) );
  AOI22X1TF U690 ( .A0(IO_DATAINB[6]), .A1(N246), .B0(D_ADDR[7]), .B1(N1171), 
        .Y(N357) );
  AOI211X1TF U691 ( .A0(N475), .A1(N245), .B0(N331), .C0(N330), .Y(N390) );
  AOI211X1TF U692 ( .A0(N841), .A1(N328), .B0(N842), .C0(N327), .Y(N329) );
  OAI22X1TF U693 ( .A0(N838), .A1(N837), .B0(N836), .B1(N201), .Y(N842) );
  OAI211X1TF U694 ( .A0(N393), .A1(N147), .B0(N1067), .C0(N1066), .Y(N464) );
  INVX2TF U695 ( .A(N355), .Y(N391) );
  OAI211X1TF U696 ( .A0(N872), .A1(N831), .B0(N788), .C0(N334), .Y(N355) );
  AOI211X1TF U697 ( .A0(N506), .A1(N865), .B0(N789), .C0(N333), .Y(N334) );
  INVX2TF U698 ( .A(N833), .Y(N840) );
  INVX2TF U699 ( .A(N779), .Y(N790) );
  OAI22X1TF U700 ( .A0(N785), .A1(N835), .B0(N867), .B1(N784), .Y(N789) );
  AOI211X1TF U701 ( .A0(REG_A[4]), .A1(N151), .B0(N781), .C0(N780), .Y(N785)
         );
  AOI22X1TF U702 ( .A0(N142), .A1(N787), .B0(REG_A[2]), .B1(N786), .Y(N788) );
  OAI21X1TF U703 ( .A0(N142), .A1(N139), .B0(N796), .Y(N786) );
  AOI22X1TF U704 ( .A0(IO_DATAINB[2]), .A1(N389), .B0(D_ADDR[3]), .B1(N173), 
        .Y(N1067) );
  INVX2TF U705 ( .A(N356), .Y(N393) );
  AOI21X1TF U706 ( .A0(N471), .A1(N245), .B0(N336), .Y(N338) );
  OAI211X1TF U707 ( .A0(N228), .A1(N774), .B0(N773), .C0(N772), .Y(N775) );
  OAI32X1TF U708 ( .A0(N200), .A1(REG_B[1]), .A2(N139), .B0(N796), .B1(N200), 
        .Y(N777) );
  INVX2TF U709 ( .A(N838), .Y(N769) );
  AOI21X1TF U710 ( .A0(IO_DATAINA[0]), .A1(N192), .B0(N379), .Y(N380) );
  OAI211X1TF U711 ( .A0(N392), .A1(N148), .B0(N378), .C0(N377), .Y(N379) );
  NOR2X1TF U712 ( .A(N42), .B(N1118), .Y(N1140) );
  AOI22X1TF U713 ( .A0(IO_DATAINB[0]), .A1(N246), .B0(D_ADDR[1]), .B1(N1171), 
        .Y(N378) );
  AND2X2TF U714 ( .A(N243), .B(N354), .Y(N389) );
  AND2X2TF U715 ( .A(N417), .B(N353), .Y(N354) );
  INVX2TF U716 ( .A(N1032), .Y(N353) );
  AOI211X1TF U717 ( .A0(REG_A[0]), .A1(N325), .B0(N324), .C0(N323), .Y(N392)
         );
  OAI211X1TF U718 ( .A0(N861), .A1(N862), .B0(N858), .C0(N322), .Y(N323) );
  AOI22X1TF U719 ( .A0(N244), .A1(N504), .B0(N470), .B1(N245), .Y(N322) );
  OAI31X1TF U720 ( .A0(N857), .A1(N856), .A2(N855), .B0(N854), .Y(N858) );
  NOR2X1TF U721 ( .A(N247), .B(N216), .Y(N855) );
  NOR2X1TF U722 ( .A(N853), .B(N200), .Y(N856) );
  NOR4BX1TF U723 ( .AN(N830), .B(N829), .C(N828), .D(N827), .Y(N846) );
  NOR2X1TF U724 ( .A(N145), .B(N228), .Y(N828) );
  OAI22X1TF U725 ( .A0(REG_A[0]), .A1(N139), .B0(N845), .B1(N213), .Y(N321) );
  OAI21X1TF U726 ( .A0(REG_B[0]), .A1(N139), .B0(N320), .Y(N325) );
  OAI211X1TF U727 ( .A0(N863), .A1(N864), .B0(N312), .C0(N311), .Y(N313) );
  NOR3X1TF U728 ( .A(N310), .B(N873), .C(N309), .Y(N311) );
  AOI22X1TF U729 ( .A0(N43), .A1(N783), .B0(N782), .B1(N140), .Y(N867) );
  OAI211X1TF U730 ( .A0(N145), .A1(N214), .B0(N748), .C0(N747), .Y(N782) );
  INVX2TF U731 ( .A(N861), .Y(N866) );
  OAI22X1TF U732 ( .A0(N872), .A1(N871), .B0(N870), .B1(N214), .Y(N873) );
  OAI211X1TF U733 ( .A0(N446), .A1(N411), .B0(N283), .C0(N282), .Y(N284) );
  AOI211X1TF U734 ( .A0(REG_A[12]), .A1(N281), .B0(N280), .C0(N279), .Y(N282)
         );
  OAI211X1TF U735 ( .A0(N218), .A1(N145), .B0(N454), .C0(N429), .Y(N848) );
  OAI211X1TF U736 ( .A0(N212), .A1(N774), .B0(N748), .C0(N816), .Y(N428) );
  NOR2X1TF U737 ( .A(N771), .B(N450), .Y(N280) );
  INVX2TF U738 ( .A(N832), .Y(N431) );
  AOI211X1TF U739 ( .A0(REG_A[4]), .A1(N422), .B0(N781), .C0(N430), .Y(N832)
         );
  OAI22X1TF U740 ( .A0(N774), .A1(N200), .B0(N247), .B1(N216), .Y(N430) );
  NOR2X1TF U741 ( .A(N853), .B(N211), .Y(N781) );
  NOR2X1TF U742 ( .A(N145), .B(N213), .Y(N820) );
  INVX2TF U743 ( .A(N821), .Y(N432) );
  NOR4X1TF U744 ( .A(N743), .B(N780), .C(N818), .D(N827), .Y(N821) );
  NOR2X1TF U745 ( .A(N233), .B(N247), .Y(N827) );
  NOR2X1TF U746 ( .A(N144), .B(N232), .Y(N818) );
  NOR2X1TF U747 ( .A(N774), .B(N201), .Y(N780) );
  NOR2X1TF U748 ( .A(N853), .B(N215), .Y(N743) );
  INVX2TF U749 ( .A(N139), .Y(N252) );
  AOI211X1TF U750 ( .A0(REG_A[13]), .A1(N275), .B0(N274), .C0(N273), .Y(N276)
         );
  OAI21X1TF U751 ( .A0(N838), .A1(N835), .B0(N272), .Y(N273) );
  AOI211X1TF U752 ( .A0(N271), .A1(N841), .B0(N270), .C0(N269), .Y(N272) );
  AOI31X1TF U753 ( .A0(N766), .A1(N754), .A2(N753), .B0(N831), .Y(N269) );
  NOR2X1TF U754 ( .A(N864), .B(N806), .Y(N270) );
  NOR4BBX1TF U755 ( .AN(N762), .BN(N767), .C(N750), .D(N791), .Y(N806) );
  NOR2X1TF U756 ( .A(N233), .B(N774), .Y(N791) );
  NOR2X1TF U757 ( .A(N232), .B(N853), .Y(N750) );
  OAI22X1TF U758 ( .A0(N140), .A1(N770), .B0(N807), .B1(N43), .Y(N841) );
  AOI211X1TF U759 ( .A0(REG_A[2]), .A1(N746), .B0(N425), .C0(N792), .Y(N807)
         );
  NOR2X1TF U760 ( .A(N853), .B(N228), .Y(N792) );
  OAI22X1TF U761 ( .A0(N145), .A1(N201), .B0(N247), .B1(N211), .Y(N425) );
  INVX2TF U762 ( .A(N803), .Y(N271) );
  AOI21X1TF U763 ( .A0(N422), .A1(REG_A[13]), .B0(N426), .Y(N838) );
  OAI22X1TF U764 ( .A0(N247), .A1(N220), .B0(N853), .B1(N202), .Y(N426) );
  NOR4BX1TF U765 ( .AN(N5040), .B(N494), .C(N499), .D(N285), .Y(N286) );
  NOR3X1TF U766 ( .A(N742), .B(REG_B[3]), .C(N861), .Y(N285) );
  AOI221X1TF U767 ( .A0(REG_B[0]), .A1(N220), .B0(N1129), .B1(N202), .C0(
        REG_B[1]), .Y(N783) );
  AOI31X1TF U768 ( .A0(N458), .A1(N815), .A2(N454), .B0(N831), .Y(N499) );
  OAI22X1TF U769 ( .A0(N490), .A1(N771), .B0(N415), .B1(N4850), .Y(N494) );
  INVX2TF U770 ( .A(N872), .Y(N4760) );
  AOI21X1TF U771 ( .A0(N422), .A1(REG_A[2]), .B0(N4710), .Y(N872) );
  OAI22X1TF U772 ( .A0(N247), .A1(N213), .B0(N853), .B1(N200), .Y(N4710) );
  NOR4X1TF U773 ( .A(N744), .B(N857), .C(N463), .D(N829), .Y(N863) );
  NOR2X1TF U774 ( .A(N853), .B(N201), .Y(N829) );
  INVX2TF U775 ( .A(N5160), .Y(N853) );
  NOR2X1TF U776 ( .A(N247), .B(N228), .Y(N463) );
  NOR2X1TF U777 ( .A(N774), .B(N211), .Y(N857) );
  NOR2X1TF U778 ( .A(N233), .B(N144), .Y(N744) );
  AOI32X1TF U779 ( .A0(N407), .A1(REG_A[14]), .A2(N415), .B0(N5090), .B1(
        REG_A[14]), .Y(N5040) );
  OAI21X1TF U780 ( .A0(N298), .A1(N220), .B0(N297), .Y(N299) );
  AOI211X1TF U781 ( .A0(N296), .A1(N758), .B0(N295), .C0(N294), .Y(N297) );
  AOI21X1TF U782 ( .A0(N293), .A1(N292), .B0(N831), .Y(N294) );
  AOI22X1TF U783 ( .A0(REG_A[14]), .A1(N5160), .B0(REG_A[13]), .B1(N151), .Y(
        N293) );
  NOR2X1TF U784 ( .A(N291), .B(N771), .Y(N295) );
  INVX2TF U785 ( .A(N398), .Y(N771) );
  NOR2X1TF U786 ( .A(N230), .B(N140), .Y(N847) );
  OAI211X1TF U787 ( .A0(N211), .A1(N145), .B0(N773), .C0(N5150), .Y(N749) );
  NOR2X2TF U788 ( .A(N43), .B(N230), .Y(N849) );
  INVX2TF U789 ( .A(N759), .Y(N332) );
  NOR4BX1TF U790 ( .AN(N765), .B(N752), .C(N5190), .D(N5170), .Y(N759) );
  NOR2X1TF U791 ( .A(N247), .B(N201), .Y(N5170) );
  NOR2X1TF U792 ( .A(N774), .B(N228), .Y(N5190) );
  INVX2TF U793 ( .A(N746), .Y(N774) );
  NOR2X1TF U794 ( .A(N145), .B(N215), .Y(N752) );
  NOR2X2TF U795 ( .A(N1129), .B(REG_B[1]), .Y(N5160) );
  NOR2X1TF U796 ( .A(N145), .B(N222), .Y(N5120) );
  NOR2X1TF U797 ( .A(N212), .B(N247), .Y(N751) );
  INVX2TF U798 ( .A(N864), .Y(N296) );
  NAND2X2TF U799 ( .A(N398), .B(N851), .Y(N864) );
  NOR2X2TF U800 ( .A(REG_B[3]), .B(N140), .Y(N851) );
  AOI21X1TF U801 ( .A0(N412), .A1(N251), .B0(N290), .Y(N298) );
  INVX2TF U802 ( .A(N320), .Y(N290) );
  INVX2TF U803 ( .A(N854), .Y(N835) );
  INVX2TF U804 ( .A(N831), .Y(N341) );
  OR2X2TF U805 ( .A(N335), .B(N43), .Y(N831) );
  AND2X2TF U806 ( .A(N1034), .B(N256), .Y(N398) );
  AND2X2TF U807 ( .A(N158), .B(N1004), .Y(N256) );
  INVX2TF U808 ( .A(N876), .Y(N1032) );
  OAI211X1TF U809 ( .A0(N882), .A1(N1033), .B0(N869), .C0(N427), .Y(N537) );
  INVX2TF U810 ( .A(N1034), .Y(N879) );
  NOR3X1TF U811 ( .A(N210), .B(N881), .C(N1007), .Y(N1017) );
  INVX2TF U812 ( .A(N1008), .Y(N881) );
  OR2X2TF U813 ( .A(N260), .B(N259), .Y(N865) );
  NOR2X1TF U814 ( .A(N741), .B(N1033), .Y(N259) );
  INVX2TF U815 ( .A(N417), .Y(N1033) );
  OR2X2TF U816 ( .A(N1011), .B(N42), .Y(N741) );
  AOI21X1TF U817 ( .A0(N258), .A1(N878), .B0(N1006), .Y(N260) );
  INVX2TF U818 ( .A(N1007), .Y(N257) );
  NAND2BX2TF U819 ( .AN(CODE_TYPE[4]), .B(CODE_TYPE[3]), .Y(N1006) );
  AOI211X1TF U820 ( .A0(CODE_TYPE[2]), .A1(N264), .B0(CODE_TYPE[3]), .C0(N263), 
        .Y(N265) );
  INVX2TF U821 ( .A(N1009), .Y(N263) );
  OAI21X1TF U822 ( .A0(N42), .A1(N219), .B0(N261), .Y(N262) );
  INVX2TF U823 ( .A(N544), .Y(N261) );
  NOR2X1TF U824 ( .A(N569), .B(N250), .Y(N544) );
  INVX2TF U825 ( .A(N552), .Y(N254) );
  OAI22X1TF U826 ( .A0(N659), .A1(N161), .B0(N159), .B1(N627), .Y(N1112) );
  OAI22X1TF U827 ( .A0(N675), .A1(N154), .B0(N152), .B1(N200), .Y(N1113) );
  OAI22X1TF U828 ( .A0(N646), .A1(N161), .B0(N160), .B1(N614), .Y(N1102) );
  OAI22X1TF U829 ( .A0(N662), .A1(N154), .B0(N153), .B1(N202), .Y(N1103) );
  OAI22X1TF U830 ( .A0(N649), .A1(N162), .B0(N160), .B1(N617), .Y(N1156) );
  OAI22X1TF U831 ( .A0(N665), .A1(N155), .B0(N153), .B1(N222), .Y(N1157) );
  OAI22X1TF U832 ( .A0(N645), .A1(N162), .B0(N160), .B1(N613), .Y(N1122) );
  OAI22X1TF U833 ( .A0(N661), .A1(N155), .B0(N153), .B1(N220), .Y(N1123) );
  OAI22X1TF U834 ( .A0(N648), .A1(N162), .B0(N159), .B1(N6160), .Y(N1145) );
  OAI22X1TF U835 ( .A0(N664), .A1(N155), .B0(N152), .B1(N218), .Y(N1146) );
  OAI22X1TF U836 ( .A0(N647), .A1(N162), .B0(N160), .B1(N615), .Y(N1068) );
  OAI22X1TF U837 ( .A0(N663), .A1(N155), .B0(N153), .B1(N217), .Y(N1069) );
  OAI22X1TF U838 ( .A0(N658), .A1(N161), .B0(N159), .B1(N626), .Y(N1060) );
  OAI22X1TF U839 ( .A0(N674), .A1(N154), .B0(N152), .B1(N216), .Y(N1061) );
  OAI22X1TF U840 ( .A0(N653), .A1(N161), .B0(N160), .B1(N621), .Y(N1167) );
  OAI22X1TF U841 ( .A0(N669), .A1(N155), .B0(N152), .B1(N215), .Y(N1168) );
  OAI22X1TF U842 ( .A0(N650), .A1(N161), .B0(N159), .B1(N618), .Y(N1084) );
  OAI22X1TF U843 ( .A0(N666), .A1(N155), .B0(N152), .B1(N214), .Y(N1085) );
  OAI22X1TF U844 ( .A0(N651), .A1(N161), .B0(N159), .B1(N619), .Y(N1074) );
  OAI22X1TF U845 ( .A0(N667), .A1(N154), .B0(N152), .B1(N212), .Y(N1075) );
  OAI22X1TF U846 ( .A0(N657), .A1(N161), .B0(N160), .B1(N625), .Y(N1094) );
  OAI22X1TF U847 ( .A0(N673), .A1(N155), .B0(N153), .B1(N211), .Y(N1095) );
  OAI22X1TF U848 ( .A0(N652), .A1(N162), .B0(N160), .B1(N620), .Y(N1050) );
  OAI22X1TF U849 ( .A0(N668), .A1(N155), .B0(N153), .B1(N232), .Y(N1051) );
  OAI22X1TF U850 ( .A0(N660), .A1(N161), .B0(N160), .B1(N628), .Y(N1134) );
  OAI22X1TF U851 ( .A0(N676), .A1(N154), .B0(N153), .B1(N213), .Y(N1135) );
  OAI22X1TF U852 ( .A0(N655), .A1(N162), .B0(N159), .B1(N623), .Y(N1026) );
  OAI22X1TF U853 ( .A0(N654), .A1(N162), .B0(N159), .B1(N622), .Y(N1037) );
  OAI22X1TF U854 ( .A0(N656), .A1(N162), .B0(N159), .B1(N624), .Y(N1043) );
  AOI21X1TF U855 ( .A0(N251), .A1(N420), .B0(N143), .Y(N342) );
  AOI21X1TF U856 ( .A0(N156), .A1(N819), .B0(N420), .Y(N822) );
  AOI21X1TF U857 ( .A0(N156), .A1(N805), .B0(N418), .Y(N813) );
  AOI21X1TF U858 ( .A0(N156), .A1(N757), .B0(N409), .Y(N760) );
  OAI31X1TF U859 ( .A0(N140), .A1(N861), .A2(N797), .B0(N157), .Y(N798) );
  AOI21X1TF U860 ( .A0(N252), .A1(N424), .B0(N143), .Y(N836) );
  AOI21X1TF U861 ( .A0(N157), .A1(N326), .B0(N424), .Y(N331) );
  AOI22X1TF U862 ( .A0(N175), .A1(REG_A[5]), .B0(N251), .B1(N201), .Y(N326) );
  AOI21X1TF U863 ( .A0(N422), .A1(N854), .B0(N143), .Y(N796) );
  AOI22X1TF U864 ( .A0(N746), .A1(REG_A[13]), .B0(N150), .B1(REG_A[12]), .Y(
        N747) );
  AOI21X1TF U865 ( .A0(N252), .A1(N408), .B0(N143), .Y(N870) );
  AOI21X1TF U866 ( .A0(N156), .A1(N308), .B0(N408), .Y(N310) );
  AOI22X1TF U867 ( .A0(N410), .A1(REG_A[10]), .B0(N251), .B1(N214), .Y(N308)
         );
  AOI22X1TF U868 ( .A0(N746), .A1(REG_A[15]), .B0(N151), .B1(REG_A[14]), .Y(
        N429) );
  AOI221X1TF U869 ( .A0(N175), .A1(REG_A[12]), .B0(N407), .B1(N218), .C0(N844), 
        .Y(N446) );
  AOI21X1TF U870 ( .A0(N157), .A1(N268), .B0(N413), .Y(N274) );
  AOI22X1TF U871 ( .A0(N175), .A1(REG_A[13]), .B0(N251), .B1(N217), .Y(N268)
         );
  AOI221X1TF U872 ( .A0(N175), .A1(REG_A[14]), .B0(N407), .B1(N202), .C0(N844), 
        .Y(N4850) );
  AOI22X1TF U873 ( .A0(N746), .A1(REG_A[0]), .B0(N150), .B1(REG_A[1]), .Y(
        N5150) );
  AOI21X1TF U874 ( .A0(N157), .A1(N289), .B0(N412), .Y(N300) );
  MXI2X1TF U875 ( .A(N373), .B(N237), .S0(N1186), .Y(N435) );
  NAND2X1TF U876 ( .A(OPER3_R3[1]), .B(N889), .Y(N1180) );
  NAND2X1TF U877 ( .A(OPER3_R3[0]), .B(N886), .Y(N1177) );
  OAI32XLTF U878 ( .A0(ZF), .A1(N210), .A2(N878), .B0(N741), .B1(N239), .Y(
        N542) );
  INVX2TF U879 ( .A(N1018), .Y(N5890) );
  INVX2TF U880 ( .A(N560), .Y(N561) );
  OAI2BB1X1TF U881 ( .A0N(N192), .A1N(IO_DATAINA[4]), .B0(N364), .Y(N455) );
  OAI2BB1X1TF U882 ( .A0N(N1172), .A1N(N361), .B0(N360), .Y(N362) );
  OAI2BB1X1TF U883 ( .A0N(N192), .A1N(IO_DATAINA[8]), .B0(N367), .Y(N459) );
  NAND2X1TF U884 ( .A(N368), .B(N1174), .Y(N369) );
  OAI2BB1X1TF U885 ( .A0N(N865), .A1N(N513), .B0(N318), .Y(N319) );
  AO21X1TF U886 ( .A0(N251), .A1(N418), .B0(N143), .Y(N317) );
  OAI2BB1X1TF U887 ( .A0N(N244), .A1N(N515), .B0(N306), .Y(N307) );
  AO21X1TF U888 ( .A0(N251), .A1(N409), .B0(N143), .Y(N305) );
  OAI2BB1X1TF U889 ( .A0N(N192), .A1N(IO_DATAINA[7]), .B0(N388), .Y(N5130) );
  AOI2BB1X1TF U890 ( .A0N(N833), .A1N(N795), .B0(N351), .Y(N352) );
  OAI2BB2XLTF U891 ( .B0(N793), .B1(N835), .A0N(N473), .A1N(N245), .Y(N349) );
  OAI2BB1X1TF U892 ( .A0N(N192), .A1N(IO_DATAINA[6]), .B0(N359), .Y(N451) );
  OAI2BB1X1TF U893 ( .A0N(N509), .A1N(N865), .B0(N329), .Y(N330) );
  AO22X1TF U894 ( .A0(N839), .A1(N840), .B0(N854), .B1(N843), .Y(N327) );
  AO22X1TF U895 ( .A0(N245), .A1(N472), .B0(N790), .B1(N840), .Y(N333) );
  OAI2BB1X1TF U896 ( .A0N(REG_B[1]), .A1N(N778), .B0(N340), .Y(N356) );
  AOI2BB1X1TF U897 ( .A0N(N776), .A1N(N861), .B0(N339), .Y(N340) );
  NAND3BX1TF U898 ( .AN(N777), .B(N338), .C(N337), .Y(N339) );
  NAND2X1TF U899 ( .A(N244), .B(N505), .Y(N337) );
  OAI2BB2XLTF U900 ( .B0(N335), .B1(N229), .A0N(N854), .A1N(N775), .Y(N336) );
  NAND4X1TF U901 ( .A(N292), .B(N766), .C(N767), .D(N768), .Y(N839) );
  NAND2X1TF U902 ( .A(N1140), .B(IO_STATUS[0]), .Y(N377) );
  OA21XLTF U903 ( .A0(N844), .A1(N321), .B0(REG_B[0]), .Y(N324) );
  OAI2BB2XLTF U904 ( .B0(N868), .B1(N867), .A0N(N874), .A1N(N341), .Y(N309) );
  NAND2X1TF U905 ( .A(N514), .B(N244), .Y(N312) );
  AO22X1TF U906 ( .A0(N341), .A1(N428), .B0(N854), .B1(N848), .Y(N279) );
  AOI222XLTF U907 ( .A0(N432), .A1(N851), .B0(N847), .B1(N820), .C0(N431), 
        .C1(N849), .Y(N450) );
  AO21X1TF U908 ( .A0(N252), .A1(N411), .B0(N5090), .Y(N281) );
  NAND2X1TF U909 ( .A(N516), .B(N244), .Y(N283) );
  OAI2BB1X1TF U910 ( .A0N(N244), .A1N(N517), .B0(N276), .Y(N277) );
  NAND2X1TF U911 ( .A(N398), .B(REG_B[3]), .Y(N803) );
  AO21X1TF U912 ( .A0(N251), .A1(N413), .B0(N5090), .Y(N275) );
  OAI2BB1X1TF U913 ( .A0N(N865), .A1N(N518), .B0(N286), .Y(N287) );
  INVX2TF U914 ( .A(N427), .Y(N278) );
  NAND2X1TF U915 ( .A(N746), .B(REG_A[12]), .Y(N292) );
  MXI2X1TF U916 ( .A(N251), .B(N175), .S0(REG_A[15]), .Y(N289) );
  NAND2X1TF U917 ( .A(N1034), .B(N42), .Y(N258) );
  NAND2BX1TF U918 ( .AN(N265), .B(N538), .Y(N266) );
  AOI2BB1X1TF U919 ( .A0N(N1034), .A1N(N262), .B0(N206), .Y(N267) );
  OAI2BB1X1TF U920 ( .A0N(N206), .A1N(N569), .B0(N254), .Y(N255) );
  CLKBUFX2TF U921 ( .A(N389), .Y(N246) );
  CLKBUFX2TF U922 ( .A(N1180), .Y(N249) );
  CLKBUFX2TF U923 ( .A(N1177), .Y(N248) );
  NAND2X1TF U924 ( .A(N5160), .B(REG_A[12]), .Y(N754) );
  NAND2X1TF U925 ( .A(N746), .B(REG_A[10]), .Y(N753) );
  OAI221XLTF U926 ( .A0(N1129), .A1(REG_A[0]), .B0(REG_B[0]), .B1(REG_A[1]), 
        .C0(N193), .Y(N770) );
  NAND2X1TF U927 ( .A(N422), .B(REG_A[9]), .Y(N767) );
  NAND2X1TF U928 ( .A(CODE_TYPE[4]), .B(N555), .Y(N1009) );
  NAND2X1TF U929 ( .A(N5160), .B(REG_A[11]), .Y(N748) );
  NAND2X1TF U930 ( .A(N5160), .B(REG_A[13]), .Y(N454) );
  OAI222X1TF U931 ( .A0(N149), .A1(N397), .B0(N147), .B1(N396), .C0(N421), 
        .C1(N243), .Y(N468) );
  NAND2X1TF U932 ( .A(N151), .B(REG_A[12]), .Y(N458) );
  NAND2X1TF U933 ( .A(N746), .B(REG_A[11]), .Y(N815) );
  NAND2X1TF U934 ( .A(N783), .B(N140), .Y(N742) );
  NAND2X1TF U935 ( .A(N422), .B(REG_A[10]), .Y(N467) );
  NAND2X1TF U936 ( .A(REG_A[9]), .B(N5160), .Y(N817) );
  NAND2X1TF U937 ( .A(N746), .B(REG_A[7]), .Y(N830) );
  NAND4X1TF U938 ( .A(N745), .B(N467), .C(N817), .D(N830), .Y(N874) );
  AOI222XLTF U939 ( .A0(N4810), .A1(N849), .B0(N874), .B1(N851), .C0(N4760), 
        .C1(N847), .Y(N490) );
  OAI222X1TF U940 ( .A0(N147), .A1(N397), .B0(N149), .B1(N395), .C0(N416), 
        .C1(N243), .Y(N4860) );
  NAND2X1TF U941 ( .A(N746), .B(REG_A[8]), .Y(N764) );
  NAND2X1TF U942 ( .A(N5160), .B(REG_A[10]), .Y(N768) );
  NAND4BBX1TF U943 ( .AN(N751), .BN(N5120), .C(N764), .D(N768), .Y(N758) );
  NAND2X1TF U944 ( .A(N5160), .B(REG_A[2]), .Y(N773) );
  NAND2X1TF U945 ( .A(REG_A[6]), .B(N5160), .Y(N765) );
  NAND3X1TF U946 ( .A(N554), .B(START), .C(N207), .Y(N728) );
  NOR4XLTF U947 ( .A(N250), .B(N1011), .C(N877), .D(N557), .Y(N167) );
  NAND2X1TF U948 ( .A(N708), .B(I_ADDR[4]), .Y(N709) );
  NAND2X1TF U949 ( .A(N713), .B(I_ADDR[6]), .Y(N718) );
  NOR2BX1TF U950 ( .AN(N727), .B(N726), .Y(N168) );
  NAND2X1TF U951 ( .A(STATE[0]), .B(N223), .Y(N723) );
  NAND2X1TF U952 ( .A(N42), .B(N569), .Y(N740) );
  NOR2BX1TF U953 ( .AN(N546), .B(N726), .Y(N545) );
  NAND2X1TF U954 ( .A(N559), .B(N546), .Y(N716) );
  AO22X1TF U955 ( .A0(D_ADDR[8]), .A1(N721), .B0(I_ADDR[8]), .B1(N714), .Y(
        N548) );
  OAI221XLTF U956 ( .A0(N42), .A1(N206), .B0(N250), .B1(N417), .C0(N569), .Y(
        N551) );
  NAND2X1TF U957 ( .A(I_ADDR[1]), .B(I_ADDR[2]), .Y(N705) );
  OAI2BB2XLTF U958 ( .B0(STATE[3]), .B1(N728), .A0N(N727), .A1N(N726), .Y(N729) );
  NAND2X1TF U959 ( .A(N236), .B(N736), .Y(N1020) );
  NAND2X1TF U960 ( .A(N206), .B(N1034), .Y(N1005) );
  NAND2X1TF U961 ( .A(N866), .B(REG_B[3]), .Y(N784) );
  NAND2X1TF U962 ( .A(N422), .B(REG_A[15]), .Y(N797) );
  NAND2X1TF U963 ( .A(N866), .B(N849), .Y(N837) );
  NAND2X1TF U964 ( .A(N398), .B(N849), .Y(N871) );
  NAND4X1TF U965 ( .A(N765), .B(N764), .C(N763), .D(N762), .Y(N843) );
  AOI222XLTF U966 ( .A0(N843), .A1(N851), .B0(N839), .B1(N849), .C0(N769), 
        .C1(N847), .Y(N776) );
  NAND2X1TF U967 ( .A(N151), .B(REG_A[3]), .Y(N772) );
  AOI2BB2X1TF U968 ( .B0(REG_A[3]), .B1(N800), .A0N(N230), .A1N(N799), .Y(N801) );
  NAND4BX1TF U969 ( .AN(N818), .B(N817), .C(N816), .D(N815), .Y(N850) );
  AOI222XLTF U970 ( .A0(N852), .A1(N851), .B0(N850), .B1(N849), .C0(N848), 
        .C1(N847), .Y(N862) );
  NAND2X1TF U971 ( .A(N1014), .B(N910), .Y(N1176) );
  AOI2BB2X1TF U972 ( .B0(IO_DATAINA[2]), .B1(N192), .A0N(N391), .A1N(N149), 
        .Y(N1066) );
  NAND3X1TF U973 ( .A(N1121), .B(N1120), .C(N1119), .Y(N491) );
  AO22X1TF U974 ( .A0(N1187), .A1(N227), .B0(N1188), .B1(I_DATAIN[4]), .Y(N523) );
endmodule


module SCPU_SRAM_8BIT_ALU_SPI_TOP_VG ( CLK, RST_N, CTRL_MODE, CTRL_BGN, CPU_BGN, 
        LOAD_N, CTRL_SI, ADC_PI, CTRL_RDY, CTRL_SO, NXT, SCLK1, SCLK2, LAT, 
        SPI_SO );
  input [1:0] CTRL_MODE;
  input [9:0] ADC_PI;
  output [1:0] NXT;
  input CLK, RST_N, CTRL_BGN, CPU_BGN, LOAD_N, CTRL_SI;
  output CTRL_RDY, CTRL_SO, SCLK1, SCLK2, LAT, SPI_SO;
  wire   CEN_AFTER_MUX, WEN_AFTER_MUX, I_CLK, I_RST_N, I_CTRL_BGN, I_CPU_BGN,
         I_LOAD_N, I_CTRL_SI, I_CTRL_SO, I_SCLK1, I_SCLK2, I_SPI_SO,
         SCPU_CTRL_SPI_CEN, \SCPU_CTRL_SPI_IO_DATAOUTB[0] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[1] , \SCPU_CTRL_SPI_IO_DATAOUTB[2] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[3] , \SCPU_CTRL_SPI_IO_DATAOUTB[4] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[5] , \SCPU_CTRL_SPI_IO_DATAOUTB[6] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[7] , \SCPU_CTRL_SPI_IO_DATAOUTB[8] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[9] , \SCPU_CTRL_SPI_IO_DATAOUTB[10] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[11] , \SCPU_CTRL_SPI_IO_DATAOUTB[12] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[0] , \SCPU_CTRL_SPI_IO_DATAOUTA[1] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[2] , \SCPU_CTRL_SPI_IO_DATAOUTA[3] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[4] , \SCPU_CTRL_SPI_IO_DATAOUTA[5] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[6] , \SCPU_CTRL_SPI_IO_DATAOUTA[7] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[8] , \SCPU_CTRL_SPI_IO_DATAOUTA[9] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[10] , \SCPU_CTRL_SPI_IO_DATAOUTA[11] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[12] , \SCPU_CTRL_SPI_IO_CONTROL[0] ,
         \SCPU_CTRL_SPI_IO_CONTROL[1] , \SCPU_CTRL_SPI_IO_CONTROL[2] ,
         \SCPU_CTRL_SPI_IO_CONTROL[3] , \SCPU_CTRL_SPI_IO_CONTROL[4] ,
         \SCPU_CTRL_SPI_IO_CONTROL[5] , \SCPU_CTRL_SPI_IO_CONTROL[6] ,
         SCPU_CTRL_SPI_D_WE, SCPU_CTRL_SPI_IS_I_ADDR, SCPU_CTRL_SPI_CCT_N57,
         SCPU_CTRL_SPI_CCT_N56, SCPU_CTRL_SPI_CCT_N55, SCPU_CTRL_SPI_CCT_N53,
         SCPU_CTRL_SPI_CCT_N52, SCPU_CTRL_SPI_CCT_N51,
         SCPU_CTRL_SPI_CCT_IS_SHIFT, \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[3] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[5] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[7] , \SCPU_CTRL_SPI_CCT_REG_BITS[1] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[2] , \SCPU_CTRL_SPI_CCT_REG_BITS[3] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[4] , \SCPU_CTRL_SPI_CCT_REG_BITS[5] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[6] , \SCPU_CTRL_SPI_CCT_REG_BITS[7] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[8] , \SCPU_CTRL_SPI_CCT_REG_BITS[9] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[10] , \SCPU_CTRL_SPI_CCT_REG_BITS[11] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[12] , \SCPU_CTRL_SPI_CCT_REG_BITS[13] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[14] , \SCPU_CTRL_SPI_CCT_REG_BITS[15] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[16] , \SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ,
         SCPU_CTRL_SPI_PUT_N110, SCPU_CTRL_SPI_PUT_N109,
         SCPU_CTRL_SPI_PUT_N108, \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] , SCPU_CTRL_SPI_PUT_N27,
         SCPU_CTRL_SPI_PUT_IS_ADDR_LEN_NZ, \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ,
         \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ,
         \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] ,
         \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[4] , \SCPU_CTRL_SPI_PUT_SPI_STATE[0] ,
         \SCPU_CTRL_SPI_PUT_SPI_STATE[1] , \SCPU_CTRL_SPI_PUT_CNT_STATE[0] ,
         \SCPU_CTRL_SPI_PUT_CNT_STATE[1] , \SCPU_CTRL_SPI_PUT_CNT_STATE[2] ,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N81, N82, N83, N84, N85, N86, N87, N88, N89, N93, N95, N103,
         N105, N161, N167, N168, N192, N193, N194, N195, N196, N197, N198,
         N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N215, N216, N217, N218, N219, N221, N222,
         N223, N224, N225, N236, N237, N238, N263, N264, N265, N266, N267,
         N268, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280,
         N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, N291,
         N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302,
         N303, N304, N305, N306, N307, N308, N309, N310, N311, N312, N313,
         N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324,
         N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335,
         N336, N337, N338, N339, N340, N341, N342, N343, N344, N345, N346,
         N347, N348, N349, N350, N351, N352, N353, N354, N355, N356, N357,
         N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N368,
         N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N401,
         N402, N403, N404, N405, N406, N407, N408, N409, N410, N411, N412,
         N413, N414, N415, N416, N417, N418, N419, N420, N421, N422, N423,
         N424;
  wire   [8:0] A_AFTER_MUX;
  wire   [7:0] D_AFTER_MUX;
  wire   [7:0] Q_FROM_SRAM;
  wire   [1:0] I_CTRL_MODE;
  wire   [9:0] I_ADC_PI;
  wire   [1:0] I_NXT;
  wire   [8:0] SCPU_CTRL_SPI_A_SPI;
  wire   [12:0] SCPU_CTRL_SPI_POUT;
  wire   [12:0] SCPU_CTRL_SPI_FOUT;
  wire   [9:0] SCPU_CTRL_SPI_IO_OFFSET;
  wire   [12:0] SCPU_CTRL_SPI_IO_DATAINA;
  wire   [0:0] SCPU_CTRL_SPI_IO_STATUS;
  wire   [7:0] SCPU_CTRL_SPI_D_DATAOUT;
  wire   [8:1] SCPU_CTRL_SPI_D_ADDR;
  wire   [8:0] SCPU_CTRL_SPI_I_ADDR;
  wire   [7:0] SCPU_CTRL_SPI_D_DATAIN;
  wire   [7:0] SCPU_CTRL_SPI_I_DATAIN;
  wire   [7:1] SCPU_CTRL_SPI_PUT_SRAM_REGS;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21;

  RA1SHD_IBM512X8 sram ( .Q(Q_FROM_SRAM), .A(A_AFTER_MUX), .D(D_AFTER_MUX), 
        .CLK(I_CLK), .CEN(CEN_AFTER_MUX), .WEN(WEN_AFTER_MUX) );
  PIC ipad_clk ( .IE(1'b1), .P(CLK), .Y(I_CLK) );
  PIC ipad_rst_n ( .IE(1'b1), .P(RST_N), .Y(I_RST_N) );
  PIC ipad_ctrl_mode0 ( .IE(1'b1), .P(CTRL_MODE[0]), .Y(I_CTRL_MODE[0]) );
  PIC ipad_ctrl_mode1 ( .IE(1'b1), .P(CTRL_MODE[1]), .Y(I_CTRL_MODE[1]) );
  PIC ipad_ctrl_bgn ( .IE(1'b1), .P(CTRL_BGN), .Y(I_CTRL_BGN) );
  PIC ipad_cpu_str ( .IE(1'b1), .P(CPU_BGN), .Y(I_CPU_BGN) );
  PIC ipad_load_n ( .IE(1'b1), .P(LOAD_N), .Y(I_LOAD_N) );
  PIC ipad_ctrl_si ( .IE(1'b1), .P(CTRL_SI), .Y(I_CTRL_SI) );
  PIC ipad_adc_pi0 ( .IE(1'b1), .P(ADC_PI[0]), .Y(I_ADC_PI[0]) );
  PIC ipad_adc_pi1 ( .IE(1'b1), .P(ADC_PI[1]), .Y(I_ADC_PI[1]) );
  PIC ipad_adc_pi2 ( .IE(1'b1), .P(ADC_PI[2]), .Y(I_ADC_PI[2]) );
  PIC ipad_adc_pi3 ( .IE(1'b1), .P(ADC_PI[3]), .Y(I_ADC_PI[3]) );
  PIC ipad_adc_pi4 ( .IE(1'b1), .P(ADC_PI[4]), .Y(I_ADC_PI[4]) );
  PIC ipad_adc_pi5 ( .IE(1'b1), .P(ADC_PI[5]), .Y(I_ADC_PI[5]) );
  PIC ipad_adc_pi6 ( .IE(1'b1), .P(ADC_PI[6]), .Y(I_ADC_PI[6]) );
  PIC ipad_adc_pi7 ( .IE(1'b1), .P(ADC_PI[7]), .Y(I_ADC_PI[7]) );
  PIC ipad_adc_pi8 ( .IE(1'b1), .P(ADC_PI[8]), .Y(I_ADC_PI[8]) );
  PIC ipad_adc_pi9 ( .IE(1'b1), .P(ADC_PI[9]), .Y(I_ADC_PI[9]) );
  POC8B opad_ctrl_rdy ( .A(N223), .P(CTRL_RDY) );
  POC8B opad_ctrl_so ( .A(I_CTRL_SO), .P(CTRL_SO) );
  POC8B opad_nxt0 ( .A(I_NXT[0]), .P(NXT[0]) );
  POC8B opad_nxt1 ( .A(I_NXT[1]), .P(NXT[1]) );
  POC8B opad_sclk1 ( .A(I_SCLK1), .P(SCLK1) );
  POC8B opad_sclk2 ( .A(I_SCLK2), .P(SCLK2) );
  POC8B opad_lat ( .A(N225), .P(LAT) );
  POC8B opad_spi_so ( .A(I_SPI_SO), .P(SPI_SO) );
  SHARE_SUPERALU_VG \scpu_ctrl_spi/ALU_01  ( .CLK(I_CLK), .RST_N(I_RST_N), .X_IN(
        {\SCPU_CTRL_SPI_IO_DATAOUTA[12] , \SCPU_CTRL_SPI_IO_DATAOUTA[11] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[10] , \SCPU_CTRL_SPI_IO_DATAOUTA[9] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[8] , \SCPU_CTRL_SPI_IO_DATAOUTA[7] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[6] , \SCPU_CTRL_SPI_IO_DATAOUTA[5] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[4] , \SCPU_CTRL_SPI_IO_DATAOUTA[3] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[2] , \SCPU_CTRL_SPI_IO_DATAOUTA[1] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[0] }), .Y_IN({
        \SCPU_CTRL_SPI_IO_DATAOUTB[12] , \SCPU_CTRL_SPI_IO_DATAOUTB[11] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[10] , \SCPU_CTRL_SPI_IO_DATAOUTB[9] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[8] , \SCPU_CTRL_SPI_IO_DATAOUTB[7] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[6] , \SCPU_CTRL_SPI_IO_DATAOUTB[5] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[4] , \SCPU_CTRL_SPI_IO_DATAOUTB[3] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[2] , \SCPU_CTRL_SPI_IO_DATAOUTB[1] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[0] }), .ALU_START(N265), .ALU_TYPE({
        \SCPU_CTRL_SPI_IO_CONTROL[4] , \SCPU_CTRL_SPI_IO_CONTROL[3] , 
        \SCPU_CTRL_SPI_IO_CONTROL[2] }), .MODE_TYPE({
        \SCPU_CTRL_SPI_IO_CONTROL[1] , \SCPU_CTRL_SPI_IO_CONTROL[0] }), 
        .OFFSET(SCPU_CTRL_SPI_IO_OFFSET), .FOUT(SCPU_CTRL_SPI_FOUT), .POUT(
        SCPU_CTRL_SPI_POUT), .ALU_IS_DONE(SCPU_CTRL_SPI_IO_STATUS[0]) );
  SERIAL_CPU_8BIT_VG \scpu_ctrl_spi/uut  ( .CLK(I_CLK), .ENABLE(1'b0), .RST_N(
        I_RST_N), .START(I_CPU_BGN), .I_DATAIN(SCPU_CTRL_SPI_I_DATAIN), 
        .D_DATAIN(SCPU_CTRL_SPI_D_DATAIN), .IS_I_ADDR(SCPU_CTRL_SPI_IS_I_ADDR), 
        .NXT(I_NXT), .I_ADDR(SCPU_CTRL_SPI_I_ADDR), .D_ADDR({
        SCPU_CTRL_SPI_D_ADDR, SYNOPSYS_UNCONNECTED__0}), .D_WE(
        SCPU_CTRL_SPI_D_WE), .D_DATAOUT(SCPU_CTRL_SPI_D_DATAOUT), .IO_STATUS({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, N224, SCPU_CTRL_SPI_IO_STATUS[0]}), .IO_CONTROL({
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, \SCPU_CTRL_SPI_IO_CONTROL[6] , 
        \SCPU_CTRL_SPI_IO_CONTROL[5] , \SCPU_CTRL_SPI_IO_CONTROL[4] , 
        \SCPU_CTRL_SPI_IO_CONTROL[3] , \SCPU_CTRL_SPI_IO_CONTROL[2] , 
        \SCPU_CTRL_SPI_IO_CONTROL[1] , \SCPU_CTRL_SPI_IO_CONTROL[0] }), 
        .IO_DATAINA({1'b0, 1'b0, 1'b0, SCPU_CTRL_SPI_IO_DATAINA}), 
        .IO_DATAINB({1'b0, 1'b0, 1'b0, SCPU_CTRL_SPI_POUT}), .IO_DATAOUTA({
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, \SCPU_CTRL_SPI_IO_DATAOUTA[12] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[11] , \SCPU_CTRL_SPI_IO_DATAOUTA[10] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[9] , \SCPU_CTRL_SPI_IO_DATAOUTA[8] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[7] , \SCPU_CTRL_SPI_IO_DATAOUTA[6] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[5] , \SCPU_CTRL_SPI_IO_DATAOUTA[4] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[3] , \SCPU_CTRL_SPI_IO_DATAOUTA[2] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[1] , \SCPU_CTRL_SPI_IO_DATAOUTA[0] }), 
        .IO_DATAOUTB({SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, \SCPU_CTRL_SPI_IO_DATAOUTB[12] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[11] , \SCPU_CTRL_SPI_IO_DATAOUTB[10] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[9] , \SCPU_CTRL_SPI_IO_DATAOUTB[8] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[7] , \SCPU_CTRL_SPI_IO_DATAOUTB[6] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[5] , \SCPU_CTRL_SPI_IO_DATAOUTB[4] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[3] , \SCPU_CTRL_SPI_IO_DATAOUTB[2] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[1] , \SCPU_CTRL_SPI_IO_DATAOUTB[0] }), 
        .IO_OFFSET({SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SCPU_CTRL_SPI_IO_OFFSET}) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[7]  ( .D(N161), .RN(
        SCPU_CTRL_SPI_CCT_N57), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[7] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[5]  ( .D(N161), .RN(
        SCPU_CTRL_SPI_CCT_N55), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[5] ), .QN(N284) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[3]  ( .D(N161), .RN(
        SCPU_CTRL_SPI_CCT_N53), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[3] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[2]  ( .D(N161), .RN(
        SCPU_CTRL_SPI_CCT_N52), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[1]  ( .D(N161), .RN(
        SCPU_CTRL_SPI_CCT_N51), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[6]  ( .D(N161), .RN(
        SCPU_CTRL_SPI_CCT_N56), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[16]  ( .D(I_CTRL_SI), .E(N267), 
        .CK(I_CLK), .Q(\SCPU_CTRL_SPI_CCT_REG_BITS[16] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[15]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[16] ), .E(N267), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[15] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[14]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[15] ), .E(N267), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[14] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[13]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[14] ), .E(N267), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[13] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[12]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[13] ), .E(N267), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[12] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[11]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[12] ), .E(N267), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[11] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[10]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[11] ), .E(N267), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[10] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[9]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[10] ), .E(N267), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[9] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[8]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[9] ), .E(N267), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[8] ) );
  DFFRX2TF \scpu_ctrl_spi/put/spi_state_reg[2]  ( .D(N215), .CK(I_CLK), .RN(
        \SCPU_CTRL_SPI_IO_CONTROL[6] ), .Q(N271), .QN(N103) );
  DFFRX2TF \scpu_ctrl_spi/put/spi_state_reg[0]  ( .D(N212), .CK(I_CLK), .RN(
        \SCPU_CTRL_SPI_IO_CONTROL[6] ), .Q(\SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), 
        .QN(N273) );
  DFFRX2TF \scpu_ctrl_spi/put/spi_state_reg[1]  ( .D(N213), .CK(I_CLK), .RN(
        \SCPU_CTRL_SPI_IO_CONTROL[6] ), .Q(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), 
        .QN(N289) );
  DFFRX2TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[3]  ( .D(N211), .CK(I_CLK), 
        .RN(\SCPU_CTRL_SPI_IO_CONTROL[6] ), .Q(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ), .QN(N287) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[2]  ( .D(N40), .CK(I_CLK), 
        .SN(N39), .RN(N38), .QN(N286) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[4]  ( .D(N46), .CK(I_CLK), 
        .SN(N45), .RN(N44), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[4] ), .QN(N280)
         );
  DFFRX2TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[0]  ( .D(N208), .CK(I_CLK), 
        .RN(N291), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .QN(N278) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[1]  ( .D(N37), .CK(I_CLK), 
        .SN(N36), .RN(N35), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ), .QN(N277)
         );
  DFFRX2TF \scpu_ctrl_spi/put/cnt_state_reg[1]  ( .D(SCPU_CTRL_SPI_PUT_N109), 
        .CK(I_CLK), .RN(N291), .Q(\SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .QN(N275)
         );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[3]  ( .D(N43), .CK(I_CLK), 
        .SN(N42), .RN(N41), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] ), .QN(N274)
         );
  DFFSX2TF \scpu_ctrl_spi/put/cnt_state_reg[0]  ( .D(SCPU_CTRL_SPI_PUT_N108), 
        .CK(I_CLK), .SN(\SCPU_CTRL_SPI_IO_CONTROL[6] ), .Q(
        \SCPU_CTRL_SPI_PUT_CNT_STATE[0] ), .QN(N272) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[7]  ( .D(N192), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[7] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[6]  ( .D(N193), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[6] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[5]  ( .D(N194), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[5] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[4]  ( .D(N195), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[4] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[3]  ( .D(N196), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[3] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[2]  ( .D(N197), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[2] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[1]  ( .D(N198), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[1] ) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[7]  ( .D(N207), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[7]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[6]  ( .D(N201), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[6]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[5]  ( .D(N202), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[5]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[4]  ( .D(N203), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[4]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[3]  ( .D(N204), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[3]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[2]  ( .D(N205), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[2]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[1]  ( .D(N206), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[1]) );
  DFFTRX1TF \scpu_ctrl_spi/cct/is_shift_reg  ( .D(N167), .RN(N168), .CK(I_CLK), 
        .QN(SCPU_CTRL_SPI_CCT_IS_SHIFT) );
  DFFQX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[4]  ( .D(N218), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[0]  ( .D(N217), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[0]  ( .D(N200), .CK(I_CLK), .Q(
        I_SPI_SO) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[0]  ( .D(N199), .CK(I_CLK), .Q(
        I_CTRL_SO) );
  DFFXLTF \scpu_ctrl_spi/cct/ctrl_state_reg[0]  ( .D(N219), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .QN(N288) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[0]  ( .D(N34), .CK(I_CLK), 
        .SN(N33), .RN(N32), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ) );
  DFFNSRX4TF \scpu_ctrl_spi/put/spi_MUX_reg  ( .D(N216), .CKN(I_CLK), .SN(1'b1), .RN(1'b1), .Q(N300), .QN(N105) );
  DFFNSRX1TF \scpu_ctrl_spi/cct/D_WE_reg  ( .D(N221), .CKN(I_CLK), .SN(1'b1), 
        .RN(1'b1), .QN(N281) );
  DFFNSRX1TF \scpu_ctrl_spi/put/sram_addr_reg[5]  ( .D(N86), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[5]), .QN(N276) );
  DFFNSRX1TF \scpu_ctrl_spi/put/sram_addr_reg[6]  ( .D(N87), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[6]), .QN(N282) );
  DFFNSRX1TF \scpu_ctrl_spi/put/sram_addr_reg[7]  ( .D(N88), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[7]), .QN(N283) );
  DFFNSRXLTF \scpu_ctrl_spi/cct/CEN_reg  ( .D(N222), .CKN(I_CLK), .SN(1'b1), 
        .RN(1'b1), .Q(SCPU_CTRL_SPI_CEN) );
  DFFNSRXLTF \scpu_ctrl_spi/put/is_addr_len_nz_reg  ( .D(SCPU_CTRL_SPI_PUT_N27), .CKN(I_CLK), .SN(1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_PUT_IS_ADDR_LEN_NZ) );
  DFFNSRXLTF \scpu_ctrl_spi/put/sram_addr_reg[8]  ( .D(N89), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[8]) );
  EDFFTRXLTF \scpu_ctrl_spi/cct/ctrl_state_reg[1]  ( .RN(I_CTRL_BGN), .D(1'b1), 
        .E(N238), .CK(I_CLK), .Q(N279), .QN(N95) );
  DFFRX1TF \scpu_ctrl_spi/put/cnt_state_reg[2]  ( .D(SCPU_CTRL_SPI_PUT_N110), 
        .CK(I_CLK), .RN(N291), .Q(\SCPU_CTRL_SPI_PUT_CNT_STATE[2] ) );
  DFFRX1TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[1]  ( .D(N209), .CK(I_CLK), 
        .RN(N291), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ) );
  DFFRX1TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[2]  ( .D(N210), .CK(I_CLK), 
        .RN(N291), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[1]  ( .D(N82), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[1]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[3]  ( .D(N84), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[3]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[2]  ( .D(N83), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[2]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[4]  ( .D(N85), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[4]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[0]  ( .D(N81), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[0]), .QN(N285) );
  NOR3BX2TF U245 ( .AN(N286), .B(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .C(
        \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ), .Y(N423) );
  CLKBUFX2TF U246 ( .A(N292), .Y(N293) );
  AND2X2TF U247 ( .A(N320), .B(N281), .Y(N321) );
  AND2X1TF U248 ( .A(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .B(SCPU_CTRL_SPI_FOUT[10]), .Y(SCPU_CTRL_SPI_IO_DATAINA[10]) );
  AND2X1TF U249 ( .A(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .B(SCPU_CTRL_SPI_FOUT[11]), .Y(SCPU_CTRL_SPI_IO_DATAINA[11]) );
  AND2X1TF U250 ( .A(N265), .B(SCPU_CTRL_SPI_FOUT[12]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[12]) );
  OAI22X1TF U251 ( .A0(SCPU_CTRL_SPI_PUT_IS_ADDR_LEN_NZ), .A1(N419), .B0(N333), 
        .B1(N271), .Y(N236) );
  AOI21X1TF U252 ( .A0(N333), .A1(N271), .B0(N236), .Y(N237) );
  AOI22X1TF U253 ( .A0(N337), .A1(N237), .B0(N103), .B1(N339), .Y(N215) );
  OA21XLTF U254 ( .A0(N268), .A1(I_CTRL_MODE[0]), .B0(N322), .Y(N238) );
  AND2X1TF U269 ( .A(N418), .B(N291), .Y(SCPU_CTRL_SPI_PUT_N27) );
  NAND2XLTF U270 ( .A(N272), .B(N275), .Y(N386) );
  NAND3X1TF U271 ( .A(SCPU_CTRL_SPI_CCT_IS_SHIFT), .B(N95), .C(N268), .Y(N93)
         );
  NOR2X4TF U272 ( .A(SCPU_CTRL_SPI_CEN), .B(N263), .Y(N320) );
  AOI22X1TF U273 ( .A0(N317), .A1(SCPU_CTRL_SPI_D_ADDR[8]), .B0(N320), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[16] ), .Y(N318) );
  AOI22X1TF U274 ( .A0(N317), .A1(SCPU_CTRL_SPI_D_ADDR[2]), .B0(N320), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[10] ), .Y(N303) );
  AOI22X1TF U275 ( .A0(N317), .A1(SCPU_CTRL_SPI_D_ADDR[3]), .B0(N320), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[11] ), .Y(N305) );
  AOI22X1TF U276 ( .A0(N317), .A1(SCPU_CTRL_SPI_D_ADDR[1]), .B0(N320), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[9] ), .Y(N301) );
  AOI22X1TF U277 ( .A0(N317), .A1(SCPU_CTRL_SPI_D_ADDR[4]), .B0(N320), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[12] ), .Y(N307) );
  AOI22X1TF U278 ( .A0(N317), .A1(SCPU_CTRL_SPI_D_ADDR[5]), .B0(N320), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[13] ), .Y(N309) );
  AOI22X1TF U279 ( .A0(N317), .A1(SCPU_CTRL_SPI_D_ADDR[7]), .B0(N320), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[15] ), .Y(N313) );
  AOI22X1TF U280 ( .A0(N317), .A1(SCPU_CTRL_SPI_D_ADDR[6]), .B0(N320), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[14] ), .Y(N311) );
  NAND2XLTF U281 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[4] ), .B(N294), .Y(N45) );
  NAND2XLTF U282 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[3] ), .B(N294), .Y(N42) );
  NAND2XLTF U283 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[2] ), .B(N294), .Y(N39) );
  NAND2BXLTF U284 ( .AN(\SCPU_CTRL_SPI_IO_DATAOUTB[3] ), .B(N292), .Y(N41) );
  NAND2BXLTF U285 ( .AN(\SCPU_CTRL_SPI_IO_DATAOUTB[4] ), .B(N292), .Y(N44) );
  NAND2BXLTF U286 ( .AN(\SCPU_CTRL_SPI_IO_DATAOUTB[0] ), .B(N292), .Y(N32) );
  OAI211XLTF U287 ( .A0(\SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .A1(N336), .B0(N337), .C0(N271), .Y(N335) );
  INVX1TF U288 ( .A(N323), .Y(N324) );
  NAND2XLTF U289 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[0] ), .B(N417), .Y(N33) );
  NAND2BXLTF U290 ( .AN(\SCPU_CTRL_SPI_IO_DATAOUTB[1] ), .B(N417), .Y(N35) );
  NAND2XLTF U291 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[1] ), .B(N417), .Y(N36) );
  NAND2BXLTF U292 ( .AN(\SCPU_CTRL_SPI_IO_DATAOUTB[2] ), .B(N417), .Y(N38) );
  NAND2XLTF U293 ( .A(N404), .B(SCPU_CTRL_SPI_A_SPI[3]), .Y(N403) );
  NAND2BX2TF U294 ( .AN(SCPU_CTRL_SPI_IS_I_ADDR), .B(N263), .Y(N374) );
  INVX2TF U295 ( .A(I_CTRL_BGN), .Y(N263) );
  NAND2XLTF U296 ( .A(SCPU_CTRL_SPI_A_SPI[0]), .B(SCPU_CTRL_SPI_A_SPI[1]), .Y(
        N410) );
  INVX2TF U297 ( .A(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .Y(N290) );
  CLKBUFX2TF U298 ( .A(\SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .Y(N268) );
  OR2X2TF U299 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ), .B(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .Y(N295) );
  INVX2TF U300 ( .A(I_CTRL_BGN), .Y(N264) );
  INVX2TF U301 ( .A(N290), .Y(N265) );
  INVX2TF U302 ( .A(N93), .Y(N266) );
  INVX2TF U303 ( .A(N93), .Y(N267) );
  NOR3X4TF U304 ( .A(I_CTRL_BGN), .B(N293), .C(N351), .Y(N360) );
  NOR3X1TF U305 ( .A(N268), .B(N279), .C(N264), .Y(N325) );
  NAND4BX2TF U306 ( .AN(N222), .B(I_CTRL_BGN), .C(SCPU_CTRL_SPI_CCT_IS_SHIFT), 
        .D(N363), .Y(N373) );
  CLKBUFX2TF U307 ( .A(\SCPU_CTRL_SPI_IO_CONTROL[6] ), .Y(N291) );
  NOR3X4TF U308 ( .A(N350), .B(N349), .C(N293), .Y(N361) );
  NAND2X1TF U309 ( .A(N424), .B(SCPU_CTRL_SPI_PUT_IS_ADDR_LEN_NZ), .Y(N414) );
  NOR2X1TF U310 ( .A(N336), .B(N352), .Y(N348) );
  NAND2X1TF U311 ( .A(I_CTRL_BGN), .B(N323), .Y(N331) );
  NOR2X1TF U312 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[3] ), .B(N296), .Y(N167)
         );
  AOI222XLTF U313 ( .A0(N361), .A1(I_SPI_SO), .B0(N360), .B1(Q_FROM_SRAM[0]), 
        .C0(SCPU_CTRL_SPI_PUT_SRAM_REGS[1]), .C1(N359), .Y(N362) );
  AOI222XLTF U314 ( .A0(N361), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[3]), .B0(N360), 
        .B1(Q_FROM_SRAM[3]), .C0(N359), .C1(SCPU_CTRL_SPI_PUT_SRAM_REGS[4]), 
        .Y(N355) );
  AOI222XLTF U315 ( .A0(N361), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[5]), .B0(N360), 
        .B1(Q_FROM_SRAM[5]), .C0(N359), .C1(SCPU_CTRL_SPI_PUT_SRAM_REGS[6]), 
        .Y(N357) );
  AOI222XLTF U316 ( .A0(N361), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[4]), .B0(N360), 
        .B1(Q_FROM_SRAM[4]), .C0(N359), .C1(SCPU_CTRL_SPI_PUT_SRAM_REGS[5]), 
        .Y(N356) );
  AOI222XLTF U317 ( .A0(N361), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[1]), .B0(N360), 
        .B1(Q_FROM_SRAM[1]), .C0(N359), .C1(SCPU_CTRL_SPI_PUT_SRAM_REGS[2]), 
        .Y(N353) );
  AOI222XLTF U318 ( .A0(N361), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[2]), .B0(N360), 
        .B1(Q_FROM_SRAM[2]), .C0(N359), .C1(SCPU_CTRL_SPI_PUT_SRAM_REGS[3]), 
        .Y(N354) );
  AOI222XLTF U319 ( .A0(N361), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[6]), .B0(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[7]), .B1(N359), .C0(N360), .C1(
        Q_FROM_SRAM[6]), .Y(N358) );
  NAND3X1TF U320 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .B(
        \SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .C(N103), .Y(N351) );
  NAND2X1TF U321 ( .A(N319), .B(N318), .Y(A_AFTER_MUX[8]) );
  NAND2X1TF U322 ( .A(N314), .B(N313), .Y(A_AFTER_MUX[7]) );
  NAND2X1TF U323 ( .A(N312), .B(N311), .Y(A_AFTER_MUX[6]) );
  NAND2X1TF U324 ( .A(N310), .B(N309), .Y(A_AFTER_MUX[5]) );
  NAND2X1TF U325 ( .A(N308), .B(N307), .Y(A_AFTER_MUX[4]) );
  NAND2X1TF U326 ( .A(N306), .B(N305), .Y(A_AFTER_MUX[3]) );
  NAND2X1TF U327 ( .A(N304), .B(N303), .Y(A_AFTER_MUX[2]) );
  NAND2X1TF U328 ( .A(N302), .B(N301), .Y(A_AFTER_MUX[1]) );
  CLKBUFX2TF U329 ( .A(N417), .Y(N292) );
  INVX2TF U330 ( .A(N291), .Y(N417) );
  AO21X1TF U331 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[3] ), .A1(N296), .B0(
        N167), .Y(SCPU_CTRL_SPI_CCT_N53) );
  NAND2X1TF U332 ( .A(N424), .B(N418), .Y(N420) );
  NOR2X1TF U333 ( .A(N350), .B(N348), .Y(N385) );
  NOR2X1TF U334 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ), .B(N297), .Y(N298)
         );
  NAND2X1TF U335 ( .A(N284), .B(N326), .Y(N297) );
  NOR2X1TF U336 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ), .B(N327), .Y(N326)
         );
  INVX2TF U337 ( .A(N331), .Y(N161) );
  NAND2X1TF U338 ( .A(N167), .B(N168), .Y(N323) );
  OR3X1TF U339 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ), .B(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ), .C(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .Y(N296) );
  NOR2X2TF U340 ( .A(N293), .B(N352), .Y(N359) );
  NAND3X1TF U341 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .B(N273), .C(N271), 
        .Y(N352) );
  OAI2BB2XLTF U342 ( .B0(N339), .B1(N414), .A0N(
        \SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .A1N(N335), .Y(N213) );
  OAI2BB1X1TF U343 ( .A0N(N320), .A1N(\SCPU_CTRL_SPI_CCT_REG_BITS[8] ), .B0(
        N299), .Y(A_AFTER_MUX[0]) );
  OAI221XLTF U344 ( .A0(N105), .A1(SCPU_CTRL_SPI_A_SPI[0]), .B0(N300), .B1(
        SCPU_CTRL_SPI_I_ADDR[0]), .C0(N264), .Y(N299) );
  AO22X1TF U345 ( .A0(N321), .A1(I_CTRL_SO), .B0(SCPU_CTRL_SPI_D_DATAOUT[0]), 
        .B1(N263), .Y(D_AFTER_MUX[0]) );
  NOR2X1TF U346 ( .A(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ), .B(N334), .Y(N336)
         );
  NAND2X1TF U347 ( .A(N268), .B(N279), .Y(N222) );
  NOR2X2TF U348 ( .A(N374), .B(N300), .Y(N317) );
  NOR2X2TF U349 ( .A(N300), .B(N382), .Y(N315) );
  NAND2X2TF U350 ( .A(SCPU_CTRL_SPI_IS_I_ADDR), .B(N263), .Y(N382) );
  NOR2X2TF U351 ( .A(I_CTRL_BGN), .B(N105), .Y(N316) );
  CLKBUFX2TF U352 ( .A(N292), .Y(N294) );
  AO21X1TF U353 ( .A0(\SCPU_CTRL_SPI_IO_DATAOUTA[6] ), .A1(N417), .B0(N396), 
        .Y(N87) );
  AO22X1TF U354 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[4]), .B0(N384), .B1(I_ADC_PI[4]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[4]) );
  AO22X1TF U355 ( .A0(N265), .A1(SCPU_CTRL_SPI_FOUT[8]), .B0(N384), .B1(
        I_ADC_PI[8]), .Y(SCPU_CTRL_SPI_IO_DATAINA[8]) );
  AO22X1TF U356 ( .A0(N265), .A1(SCPU_CTRL_SPI_FOUT[9]), .B0(N384), .B1(
        I_ADC_PI[9]), .Y(SCPU_CTRL_SPI_IO_DATAINA[9]) );
  AO22X1TF U357 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[7]), .B0(N384), .B1(I_ADC_PI[7]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[7]) );
  AO22X1TF U358 ( .A0(N265), .A1(SCPU_CTRL_SPI_FOUT[6]), .B0(N384), .B1(
        I_ADC_PI[6]), .Y(SCPU_CTRL_SPI_IO_DATAINA[6]) );
  INVX2TF U359 ( .A(N265), .Y(N384) );
  AOI31X1TF U360 ( .A0(N424), .A1(N423), .A2(N274), .B0(N280), .Y(N46) );
  NOR2X1TF U361 ( .A(\SCPU_CTRL_SPI_PUT_CNT_STATE[0] ), .B(N388), .Y(
        SCPU_CTRL_SPI_PUT_N108) );
  OAI32X1TF U362 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ), .A1(
        \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .A2(N420), .B0(N421), .B1(N277), 
        .Y(N37) );
  AOI32X1TF U363 ( .A0(N424), .A1(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] ), .A2(
        N423), .B0(N422), .B1(N274), .Y(N43) );
  AOI32X1TF U364 ( .A0(N421), .A1(N422), .A2(N277), .B0(N286), .B1(N422), .Y(
        N40) );
  OAI211X1TF U365 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] ), .A1(
        \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[4] ), .B0(N424), .C0(N423), .Y(N422)
         );
  NOR2X1TF U366 ( .A(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .B(N419), .Y(N421)
         );
  OAI211X1TF U367 ( .A0(N348), .A1(N278), .B0(N351), .C0(N347), .Y(N208) );
  OAI211X1TF U368 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .A1(N347), .B0(
        N351), .C0(N346), .Y(N209) );
  OAI21X1TF U369 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .A1(N385), .B0(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .Y(N346) );
  OAI31X1TF U370 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .A1(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .A2(N385), .B0(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ), .Y(N345) );
  AOI22X1TF U371 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ), .A1(N343), .B0(
        N344), .B1(N287), .Y(N211) );
  AOI21X1TF U372 ( .A0(N349), .A1(N334), .B0(N385), .Y(N343) );
  INVX2TF U373 ( .A(N385), .Y(N387) );
  OAI21X1TF U374 ( .A0(N326), .A1(N284), .B0(N297), .Y(SCPU_CTRL_SPI_CCT_N55)
         );
  OAI22X1TF U375 ( .A0(I_CTRL_MODE[0]), .A1(N329), .B0(N328), .B1(N331), .Y(
        N218) );
  AOI21X1TF U376 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ), .A1(N327), .B0(
        N326), .Y(N328) );
  INVX2TF U377 ( .A(N167), .Y(N327) );
  OAI21X1TF U378 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .A1(N331), .B0(
        N330), .Y(N217) );
  NOR4X1TF U379 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[7] ), .B(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ), .C(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[5] ), .D(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ), .Y(N168) );
  INVX2TF U380 ( .A(N362), .Y(N200) );
  INVX2TF U381 ( .A(N355), .Y(N204) );
  INVX2TF U382 ( .A(N357), .Y(N202) );
  INVX2TF U383 ( .A(N356), .Y(N203) );
  INVX2TF U384 ( .A(N353), .Y(N206) );
  INVX2TF U385 ( .A(N354), .Y(N205) );
  INVX2TF U386 ( .A(N358), .Y(N201) );
  INVX2TF U387 ( .A(N352), .Y(N349) );
  INVX2TF U388 ( .A(N351), .Y(N350) );
  OAI21X1TF U389 ( .A0(N383), .A1(N373), .B0(N372), .Y(N192) );
  AOI22X1TF U390 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[8] ), .A1(N266), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[7] ), .B1(N371), .Y(N372) );
  OAI21X1TF U391 ( .A0(N376), .A1(N373), .B0(N365), .Y(N198) );
  AOI22X1TF U392 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[2] ), .A1(N266), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[1] ), .B1(N371), .Y(N365) );
  OAI21X1TF U393 ( .A0(N377), .A1(N373), .B0(N366), .Y(N197) );
  AOI22X1TF U394 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[3] ), .A1(N266), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[2] ), .B1(N371), .Y(N366) );
  OAI21X1TF U395 ( .A0(N378), .A1(N373), .B0(N367), .Y(N196) );
  AOI22X1TF U396 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[4] ), .A1(N266), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[3] ), .B1(N371), .Y(N367) );
  OAI21X1TF U397 ( .A0(N379), .A1(N373), .B0(N368), .Y(N195) );
  AOI22X1TF U398 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[5] ), .A1(N266), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[4] ), .B1(N371), .Y(N368) );
  OAI21X1TF U399 ( .A0(N375), .A1(N373), .B0(N364), .Y(N199) );
  AOI22X1TF U400 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[1] ), .A1(N266), .B0(
        I_CTRL_SO), .B1(N371), .Y(N364) );
  OAI21X1TF U401 ( .A0(N381), .A1(N373), .B0(N370), .Y(N193) );
  AOI22X1TF U402 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[7] ), .A1(N266), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[6] ), .B1(N371), .Y(N370) );
  OAI21X1TF U403 ( .A0(N380), .A1(N373), .B0(N369), .Y(N194) );
  AOI22X1TF U404 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[6] ), .A1(N266), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[5] ), .B1(N371), .Y(N369) );
  OAI211X4TF U405 ( .A0(N95), .A1(N363), .B0(N268), .C0(
        SCPU_CTRL_SPI_CCT_IS_SHIFT), .Y(N371) );
  INVX2TF U406 ( .A(I_CTRL_MODE[1]), .Y(N363) );
  AND2X2TF U407 ( .A(N338), .B(N271), .Y(N225) );
  NOR2X1TF U408 ( .A(N95), .B(N268), .Y(N223) );
  AND2X2TF U409 ( .A(SCPU_CTRL_SPI_CEN), .B(I_CTRL_BGN), .Y(CEN_AFTER_MUX) );
  AOI32X1TF U410 ( .A0(N105), .A1(N264), .A2(SCPU_CTRL_SPI_D_WE), .B0(
        I_CTRL_BGN), .B1(N281), .Y(WEN_AFTER_MUX) );
  NOR2X1TF U411 ( .A(N379), .B(N382), .Y(SCPU_CTRL_SPI_I_DATAIN[4]) );
  NOR2X1TF U412 ( .A(N377), .B(N382), .Y(SCPU_CTRL_SPI_I_DATAIN[2]) );
  NOR2X1TF U413 ( .A(N381), .B(N382), .Y(SCPU_CTRL_SPI_I_DATAIN[6]) );
  NOR2X1TF U414 ( .A(N376), .B(N382), .Y(SCPU_CTRL_SPI_I_DATAIN[1]) );
  NOR2X1TF U415 ( .A(N380), .B(N382), .Y(SCPU_CTRL_SPI_I_DATAIN[5]) );
  NOR2X1TF U416 ( .A(N375), .B(N382), .Y(SCPU_CTRL_SPI_I_DATAIN[0]) );
  NOR2X1TF U417 ( .A(N383), .B(N382), .Y(SCPU_CTRL_SPI_I_DATAIN[7]) );
  NOR2X1TF U418 ( .A(N378), .B(N382), .Y(SCPU_CTRL_SPI_I_DATAIN[3]) );
  NOR2X1TF U419 ( .A(N381), .B(N374), .Y(SCPU_CTRL_SPI_D_DATAIN[6]) );
  INVX2TF U420 ( .A(Q_FROM_SRAM[6]), .Y(N381) );
  NOR2X1TF U421 ( .A(N380), .B(N374), .Y(SCPU_CTRL_SPI_D_DATAIN[5]) );
  INVX2TF U422 ( .A(Q_FROM_SRAM[5]), .Y(N380) );
  NOR2X1TF U423 ( .A(N383), .B(N374), .Y(SCPU_CTRL_SPI_D_DATAIN[7]) );
  INVX2TF U424 ( .A(Q_FROM_SRAM[7]), .Y(N383) );
  NOR2X1TF U425 ( .A(N377), .B(N374), .Y(SCPU_CTRL_SPI_D_DATAIN[2]) );
  INVX2TF U426 ( .A(Q_FROM_SRAM[2]), .Y(N377) );
  NOR2X1TF U427 ( .A(N378), .B(N374), .Y(SCPU_CTRL_SPI_D_DATAIN[3]) );
  INVX2TF U428 ( .A(Q_FROM_SRAM[3]), .Y(N378) );
  NOR2X1TF U429 ( .A(N375), .B(N374), .Y(SCPU_CTRL_SPI_D_DATAIN[0]) );
  INVX2TF U430 ( .A(Q_FROM_SRAM[0]), .Y(N375) );
  NOR2X1TF U431 ( .A(N379), .B(N374), .Y(SCPU_CTRL_SPI_D_DATAIN[4]) );
  INVX2TF U432 ( .A(Q_FROM_SRAM[4]), .Y(N379) );
  NOR2X1TF U433 ( .A(N376), .B(N374), .Y(SCPU_CTRL_SPI_D_DATAIN[1]) );
  INVX2TF U434 ( .A(Q_FROM_SRAM[1]), .Y(N376) );
  OAI32X1TF U435 ( .A0(N293), .A1(N105), .A2(N332), .B0(N419), .B1(N293), .Y(
        N216) );
  INVX2TF U436 ( .A(N424), .Y(N419) );
  OAI21X1TF U437 ( .A0(N103), .A1(N341), .B0(N340), .Y(N212) );
  OAI32X1TF U438 ( .A0(N339), .A1(N411), .A2(N338), .B0(
        \SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .B1(N337), .Y(N340) );
  NOR2X1TF U439 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .B(
        \SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .Y(N338) );
  AOI21X1TF U440 ( .A0(N336), .A1(N337), .B0(\SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), 
        .Y(N341) );
  INVX2TF U441 ( .A(N339), .Y(N337) );
  AOI21X1TF U442 ( .A0(N271), .A1(N333), .B0(N388), .Y(N339) );
  NOR3X1TF U443 ( .A(\SCPU_CTRL_SPI_PUT_CNT_STATE[0] ), .B(
        \SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .C(\SCPU_CTRL_SPI_PUT_CNT_STATE[2] ), .Y(N388) );
  INVX2TF U444 ( .A(N342), .Y(N334) );
  NOR3X1TF U445 ( .A(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ), .B(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .C(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .Y(N342) );
  AOI22X1TF U446 ( .A0(SCPU_CTRL_SPI_A_SPI[8]), .A1(N316), .B0(N315), .B1(
        SCPU_CTRL_SPI_I_ADDR[8]), .Y(N319) );
  AOI22X1TF U447 ( .A0(SCPU_CTRL_SPI_A_SPI[7]), .A1(N316), .B0(N315), .B1(
        SCPU_CTRL_SPI_I_ADDR[7]), .Y(N314) );
  AOI22X1TF U448 ( .A0(SCPU_CTRL_SPI_A_SPI[6]), .A1(N316), .B0(N315), .B1(
        SCPU_CTRL_SPI_I_ADDR[6]), .Y(N312) );
  AOI22X1TF U449 ( .A0(SCPU_CTRL_SPI_A_SPI[5]), .A1(N316), .B0(N315), .B1(
        SCPU_CTRL_SPI_I_ADDR[5]), .Y(N310) );
  AOI22X1TF U450 ( .A0(SCPU_CTRL_SPI_A_SPI[4]), .A1(N316), .B0(N315), .B1(
        SCPU_CTRL_SPI_I_ADDR[4]), .Y(N308) );
  AOI22X1TF U451 ( .A0(SCPU_CTRL_SPI_A_SPI[3]), .A1(N316), .B0(N315), .B1(
        SCPU_CTRL_SPI_I_ADDR[3]), .Y(N306) );
  AOI22X1TF U452 ( .A0(SCPU_CTRL_SPI_A_SPI[2]), .A1(N316), .B0(N315), .B1(
        SCPU_CTRL_SPI_I_ADDR[2]), .Y(N304) );
  AOI22X1TF U453 ( .A0(SCPU_CTRL_SPI_A_SPI[1]), .A1(N316), .B0(N315), .B1(
        SCPU_CTRL_SPI_I_ADDR[1]), .Y(N302) );
  OAI31X1TF U454 ( .A0(SCPU_CTRL_SPI_A_SPI[3]), .A1(N416), .A2(N407), .B0(N406), .Y(N84) );
  AOI22X1TF U455 ( .A0(SCPU_CTRL_SPI_A_SPI[3]), .A1(N405), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[3] ), .B1(N294), .Y(N406) );
  AOI21X1TF U456 ( .A0(N411), .A1(N404), .B0(N294), .Y(N405) );
  OAI31X1TF U457 ( .A0(SCPU_CTRL_SPI_A_SPI[2]), .A1(N416), .A2(N410), .B0(N409), .Y(N83) );
  AOI22X1TF U458 ( .A0(SCPU_CTRL_SPI_A_SPI[2]), .A1(N408), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[2] ), .B1(N293), .Y(N409) );
  AOI31X1TF U459 ( .A0(N411), .A1(SCPU_CTRL_SPI_A_SPI[0]), .A2(
        SCPU_CTRL_SPI_A_SPI[1]), .B0(N294), .Y(N408) );
  OAI31X1TF U460 ( .A0(SCPU_CTRL_SPI_A_SPI[1]), .A1(N416), .A2(N285), .B0(N413), .Y(N82) );
  AOI22X1TF U461 ( .A0(SCPU_CTRL_SPI_A_SPI[1]), .A1(N412), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[1] ), .B1(N293), .Y(N413) );
  AOI21X1TF U462 ( .A0(N411), .A1(SCPU_CTRL_SPI_A_SPI[0]), .B0(N294), .Y(N412)
         );
  OAI31X1TF U463 ( .A0(SCPU_CTRL_SPI_A_SPI[4]), .A1(N416), .A2(N403), .B0(N402), .Y(N85) );
  AOI22X1TF U464 ( .A0(SCPU_CTRL_SPI_A_SPI[4]), .A1(N401), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[4] ), .B1(N294), .Y(N402) );
  AOI31X1TF U465 ( .A0(N411), .A1(N404), .A2(SCPU_CTRL_SPI_A_SPI[3]), .B0(N294), .Y(N401) );
  OAI21X1TF U466 ( .A0(SCPU_CTRL_SPI_A_SPI[0]), .A1(N416), .B0(N415), .Y(N81)
         );
  AOI32X1TF U467 ( .A0(SCPU_CTRL_SPI_A_SPI[0]), .A1(N291), .A2(N414), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[0] ), .B1(N293), .Y(N415) );
  OAI21X1TF U468 ( .A0(SCPU_CTRL_SPI_A_SPI[5]), .A1(N400), .B0(N399), .Y(N86)
         );
  AOI22X1TF U469 ( .A0(SCPU_CTRL_SPI_A_SPI[5]), .A1(N398), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[5] ), .B1(N294), .Y(N399) );
  OAI31X1TF U470 ( .A0(SCPU_CTRL_SPI_A_SPI[8]), .A1(N283), .A2(N392), .B0(N391), .Y(N89) );
  AOI22X1TF U471 ( .A0(SCPU_CTRL_SPI_A_SPI[8]), .A1(N390), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[8] ), .B1(N293), .Y(N391) );
  OAI21X1TF U472 ( .A0(SCPU_CTRL_SPI_A_SPI[7]), .A1(N416), .B0(N394), .Y(N390)
         );
  OAI21X1TF U473 ( .A0(N394), .A1(N283), .B0(N393), .Y(N88) );
  NOR3X1TF U474 ( .A(N397), .B(N276), .C(N282), .Y(N389) );
  OAI32X1TF U475 ( .A0(SCPU_CTRL_SPI_A_SPI[6]), .A1(N276), .A2(N400), .B0(N395), .B1(N282), .Y(N396) );
  OAI31X1TF U476 ( .A0(N414), .A1(N397), .A2(N276), .B0(N291), .Y(N395) );
  OR2X2TF U477 ( .A(N397), .B(N416), .Y(N400) );
  NAND2X2TF U478 ( .A(N291), .B(N411), .Y(N416) );
  INVX2TF U479 ( .A(N414), .Y(N411) );
  AND3X2TF U480 ( .A(N289), .B(\SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .C(N103), 
        .Y(N424) );
  INVX2TF U481 ( .A(N407), .Y(N404) );
  AND2X2TF U482 ( .A(N332), .B(N271), .Y(N224) );
  NOR2X1TF U483 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .B(N273), .Y(N332) );
  NOR3X1TF U484 ( .A(N105), .B(N275), .C(N272), .Y(I_SCLK1) );
  NOR3X1TF U485 ( .A(\SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .B(N105), .C(N272), 
        .Y(I_SCLK2) );
  OAI2BB1X1TF U486 ( .A0N(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .A1N(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ), .B0(N295), .Y(
        SCPU_CTRL_SPI_CCT_N51) );
  OAI2BB1X1TF U487 ( .A0N(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ), .A1N(N295), 
        .B0(N296), .Y(SCPU_CTRL_SPI_CCT_N52) );
  AO21X1TF U488 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ), .A1(N297), .B0(
        N298), .Y(SCPU_CTRL_SPI_CCT_N56) );
  XOR2X1TF U489 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[7] ), .B(N298), .Y(
        SCPU_CTRL_SPI_CCT_N57) );
  AO22X1TF U490 ( .A0(N321), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[1] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[1]), .B1(N264), .Y(D_AFTER_MUX[1]) );
  AO22X1TF U491 ( .A0(N321), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[2] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[2]), .B1(N264), .Y(D_AFTER_MUX[2]) );
  AO22X1TF U492 ( .A0(N321), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[3] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[3]), .B1(N264), .Y(D_AFTER_MUX[3]) );
  AO22X1TF U493 ( .A0(N321), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[4] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[4]), .B1(N264), .Y(D_AFTER_MUX[4]) );
  AO22X1TF U494 ( .A0(N321), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[5] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[5]), .B1(N264), .Y(D_AFTER_MUX[5]) );
  AO22X1TF U495 ( .A0(N321), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[6] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[6]), .B1(N264), .Y(D_AFTER_MUX[6]) );
  AO22X1TF U496 ( .A0(N321), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[7] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[7]), .B1(N264), .Y(D_AFTER_MUX[7]) );
  NAND2BX1TF U497 ( .AN(N222), .B(I_CTRL_MODE[1]), .Y(N221) );
  OAI221XLTF U498 ( .A0(N268), .A1(I_LOAD_N), .B0(N288), .B1(N323), .C0(
        I_CTRL_BGN), .Y(N322) );
  AO22X1TF U499 ( .A0(N268), .A1(N161), .B0(N325), .B1(N322), .Y(N219) );
  NAND3BX1TF U500 ( .AN(I_LOAD_N), .B(N325), .C(N324), .Y(N329) );
  AO21X1TF U501 ( .A0(I_CTRL_MODE[0]), .A1(I_CTRL_MODE[1]), .B0(N329), .Y(N330) );
  NAND2X1TF U502 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .B(N273), .Y(N333) );
  NAND2X1TF U503 ( .A(N342), .B(N348), .Y(N344) );
  NAND3X1TF U504 ( .A(N351), .B(N345), .C(N344), .Y(N210) );
  NAND2X1TF U505 ( .A(N348), .B(N278), .Y(N347) );
  AO22X1TF U506 ( .A0(N361), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[7]), .B0(
        Q_FROM_SRAM[7]), .B1(N360), .Y(N207) );
  AO22X1TF U507 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[0]), .B0(N384), .B1(I_ADC_PI[0]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[0]) );
  AO22X1TF U508 ( .A0(N265), .A1(SCPU_CTRL_SPI_FOUT[1]), .B0(N384), .B1(
        I_ADC_PI[1]), .Y(SCPU_CTRL_SPI_IO_DATAINA[1]) );
  AO22X1TF U509 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[2]), .B0(N384), .B1(I_ADC_PI[2]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[2]) );
  AO22X1TF U510 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[3]), .B0(N384), .B1(I_ADC_PI[3]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[3]) );
  AO22X1TF U511 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[5]), .B0(N384), .B1(I_ADC_PI[5]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[5]) );
  AO22X1TF U512 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .A1(
        \SCPU_CTRL_SPI_PUT_CNT_STATE[0] ), .B0(N275), .B1(
        SCPU_CTRL_SPI_PUT_N108), .Y(SCPU_CTRL_SPI_PUT_N109) );
  AO22X1TF U513 ( .A0(N388), .A1(N387), .B0(\SCPU_CTRL_SPI_PUT_CNT_STATE[2] ), 
        .B1(N386), .Y(SCPU_CTRL_SPI_PUT_N110) );
  NAND3X1TF U514 ( .A(N280), .B(N274), .C(N423), .Y(N418) );
  NAND3X1TF U515 ( .A(SCPU_CTRL_SPI_A_SPI[2]), .B(SCPU_CTRL_SPI_A_SPI[0]), .C(
        SCPU_CTRL_SPI_A_SPI[1]), .Y(N407) );
  NAND3X1TF U516 ( .A(SCPU_CTRL_SPI_A_SPI[4]), .B(N404), .C(
        SCPU_CTRL_SPI_A_SPI[3]), .Y(N397) );
  NAND2BX1TF U517 ( .AN(N416), .B(N389), .Y(N392) );
  AO21X1TF U518 ( .A0(N411), .A1(N389), .B0(N417), .Y(N394) );
  AOI2BB2X1TF U519 ( .B0(\SCPU_CTRL_SPI_IO_DATAOUTA[7] ), .B1(N293), .A0N(
        SCPU_CTRL_SPI_A_SPI[7]), .A1N(N392), .Y(N393) );
  AOI2BB1X1TF U520 ( .A0N(N414), .A1N(N397), .B0(N292), .Y(N398) );
  XNOR2X1TF U522 ( .A(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .B(N420), .Y(N34)
         );
endmodule

