
module SHARE_SUPERALU_VG ( CLK, RST_N, X_IN, Y_IN, ALU_START, ALU_TYPE, MODE_TYPE, 
        OFFSET, FOUT, POUT, ALU_IS_DONE );
  input [12:0] X_IN;
  input [12:0] Y_IN;
  input [2:0] ALU_TYPE;
  input [1:0] MODE_TYPE;
  input [9:0] OFFSET;
  output [12:0] FOUT;
  output [12:0] POUT;
  input CLK, RST_N, ALU_START;
  output ALU_IS_DONE;
  wire   POST_WORK, PRE_WORK, \INDEX[2] , \RSHT_BITS[3] , SIGN_Y, C152_DATA4_0,
         C152_DATA4_1, C152_DATA4_2, C152_DATA4_3, C152_DATA4_4, C152_DATA4_5,
         C152_DATA4_6, C152_DATA4_7, C152_DATA4_8, C152_DATA4_9, C152_DATA4_10,
         C152_DATA4_11, N73, N74, N90, N91, N92, N121, N122, N123, N124, N128,
         N129, N657, N658, N659, N660, N661, N662, N663, N664, N665, N666,
         N667, N668, N669, N670, N671, N672, N673, N674, N675, N676, N677,
         N678, N679, N680, N681, N682, N683, N684, N685, N686, N687, N688,
         N689, N690, N691, N692, N693, N694, N695, N696, N697, N698, N699,
         N700, N701, N702, N703, N704, N705, N706, N707, N708, N709, N710,
         N711, N712, N713, N714, N715, N716, N717, N718, N719, N720, N721,
         N722, N723, N724, N725, N726, C2_Z_11, C2_Z_10, C2_Z_9, C2_Z_8,
         C2_Z_7, C2_Z_6, C2_Z_5, C2_Z_4, C2_Z_3, C2_Z_2, C2_Z_1, C2_Z_0,
         DP_OP_333_124_4748_N57, DP_OP_333_124_4748_N43,
         DP_OP_333_124_4748_N29, DP_OP_333_124_4748_N28,
         DP_OP_333_124_4748_N27, DP_OP_333_124_4748_N26,
         DP_OP_333_124_4748_N25, DP_OP_333_124_4748_N24,
         DP_OP_333_124_4748_N23, DP_OP_333_124_4748_N22,
         DP_OP_333_124_4748_N21, DP_OP_333_124_4748_N20,
         DP_OP_333_124_4748_N19, DP_OP_333_124_4748_N18,
         DP_OP_333_124_4748_N12, DP_OP_333_124_4748_N11,
         DP_OP_333_124_4748_N10, DP_OP_333_124_4748_N9, DP_OP_333_124_4748_N8,
         DP_OP_333_124_4748_N7, DP_OP_333_124_4748_N6, DP_OP_333_124_4748_N5,
         DP_OP_333_124_4748_N4, DP_OP_333_124_4748_N3, DP_OP_333_124_4748_N2,
         DP_OP_333_124_4748_N1, INTADD_0_CI, \INTADD_0_SUM[6] ,
         \INTADD_0_SUM[5] , \INTADD_0_SUM[4] , \INTADD_0_SUM[3] ,
         \INTADD_0_SUM[2] , \INTADD_0_SUM[1] , \INTADD_0_SUM[0] , INTADD_0_N7,
         INTADD_0_N6, INTADD_0_N5, INTADD_0_N4, INTADD_0_N3, INTADD_0_N2,
         INTADD_0_N1, ADD_X_132_1_N13, ADD_X_132_1_N12, ADD_X_132_1_N11,
         ADD_X_132_1_N10, ADD_X_132_1_N9, ADD_X_132_1_N8, ADD_X_132_1_N7,
         ADD_X_132_1_N6, ADD_X_132_1_N5, ADD_X_132_1_N4, ADD_X_132_1_N3,
         ADD_X_132_1_N2, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12,
         N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26,
         N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40,
         N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54,
         N55, N56, N58, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104,
         N105, N106, N107, N108, N109, N110, N111, N112, N113, N114, N115,
         N116, N117, N118, N119, N120, N125, N126, N127, N130, N131, N132,
         N133, N134, N135, N136, N137, N138, N139, N140, N141, N142, N143,
         N144, N145, N146, N147, N148, N149, N150, N151, N152, N153, N154,
         N155, N156, N157, N158, N159, N160, N161, N162, N163, N164, N165,
         N166, N167, N168, N169, N170, N171, N172, N173, N174, N175, N176,
         N177, N178, N179, N180, N181, N182, N183, N184, N185, N186, N187,
         N188, N189, N190, N191, N192, N193, N194, N195, N196, N197, N198,
         N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N214, N215, N216, N217, N218, N219, N220,
         N221, N222, N223, N224, N225, N226, N227, N228, N229, N230, N231,
         N232, N233, N234, N235, N236, N237, N238, N239, N240, N241, N242,
         N243, N244, N245, N246, N247, N248, N249, N250, N251, N252, N253,
         N254, N255, N256, N257, N258, N259, N260, N261, N262, N263, N264,
         N265, N266, N267, N268, N269, N270, N271, N272, N273, N274, N275,
         N276, N277, N278, N279, N280, N281, N282, N283, N284, N285, N286,
         N287, N288, N289, N290, N291, N292, N293, N294, N295, N296, N297,
         N298, N299, N300, N301, N302, N303, N304, N305, N306, N307, N308,
         N309, N310, N311, N312, N313, N314, N315, N316, N317, N318, N319,
         N320, N321, N322, N323, N324, N325, N326, N327, N328, N329, N330,
         N331, N332, N333, N334, N335, N336, N337, N338, N339, N340, N341,
         N342, N343, N344, N345, N346, N347, N348, N349, N350, N351, N352,
         N353, N354, N355, N356, N357, N358, N359, N360, N361, N362, N363,
         N364, N365, N366, N367, N368, N369, N370, N371, N372, N373, N374,
         N375, N376, N377, N378, N379, N380, N381, N382, N383, N384, N385,
         N386, N387, N388, N389, N390, N391, N392, N393, N394, N395, N396,
         N397, N398, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N408, N409, N410, N411, N412, N413, N414, N415, N416, N417, N418,
         N419, N420, N421, N422, N423, N424, N425, N426, N427, N428, N429,
         N430, N431, N432, N433, N434, N435, N436, N437, N438, N439, N440,
         N441, N442, N443, N444, N445, N446, N447, N448, N449, N450, N451,
         N452, N453, N454, N455, N456, N457, N458, N459, N460, N461, N462,
         N463, N464, N465, N466, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N487, N488, N489, N490, N491, N492, N493, N494, N495,
         N496, N497, N498, N499, N500, N501, N502, N503, N504, N505, N506,
         N507, N508, N509, N510, N511, N512, N513, N514, N515, N516, N517,
         N518, N519, N520, N521, N522, N523, N524, N525, N526, N527, N528,
         N529, N530, N531, N532, N533, N534, N535, N536, N537, N538, N539,
         N540, N541, N542, N543, N544, N545, N546, N547, N548, N549, N550,
         N551, N552, N553, N554, N555, N556, N557, N558, N559, N560, N561,
         N562, N563, N564, N565, N566, N567, N568, N569, N570, N571, N572,
         N573, N574, N575, N576, N577, N578, N579, N580, N581, N582, N583,
         N584, N585, N586, N587, N588, N589, N590, N591, N592, N593, N594,
         N595, N596, N597, N598, N599, N600, N601, N602, N603, N604, N605,
         N606, N607, N608, N609, N610, N611, N612, N613, N614, N615, N616,
         N617, N618, N619, N620, N621, N622, N623, N624, N625, N626, N627,
         N628, N629, N630, N631, N632, N633, N634, N635, N636, N637, N638,
         N639, N640, N641, N642, N643, N644, N645, N646, N647, N648, N649,
         N650, N651, N652, N653, N654, N655, N656, N727, N728, N729, N730,
         N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741,
         N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752,
         N753, N754, N755, N756, N757, N758, N759, N760, N761, N762, N763,
         N764, N765, N766, N767, N768, N769, N770, N771, N772, N773, N774,
         N775, N776, N777, N778, N779, N780, N781, N782, N783, N784, N785,
         N786, N787, N788, N789, N790, N791, N792, N793, N794, N795, N796,
         N797, N798, N799, N800, N801, N802, N803, N804, N805, N806, N807,
         N808, N809, N810, N811, N812, N813, N814, N815, N816, N817, N818,
         N819, N820, N821, N822, N823, N824, N825, N826, N827, N828, N829,
         N830, N831, N832, N833, N834, N835, N836, N837, N838, N839, N840,
         N841, N842, N843, N844, N845, N846, N847, N848, N849, N850, N851,
         N852, N853, N854, N855, N856, N857, N858, N859, N860, N861, N862,
         N863, N864, N865, N866, N867, N868, N869, N870, N871, N872, N873,
         N874, N875, N876, N877, N878, N879, N880, N881, N882, N883, N884,
         N885, N886, N887, N888, N889, N890, N891, N892, N893, N894, N895,
         N896, N897, N898, N899, N900, N901, N902, N903, N904, N905, N906,
         N907, N908, N909, N910, N911, N912, N913, N914, N915, N916, N917,
         N918, N919, N920, N921, N922, N923, N924, N925, N926, N927, N928,
         N929, N930, N931, N932, N933, N934, N935, N936, N937, N938, N939,
         N940, N941, N942, N943, N944, N945, N946, N947, N948, N949, N950,
         N951, N952, N953, N954, N955, N956, N957, N958, N959, N960, N961,
         N962, N963, N964, N965, N966, N967, N968, N969, N970, N971, N972,
         N973, N974, N975, N976, N977, N978, N979, N980, N981, N982, N983,
         N984, N985, N986, N987, N988, N989, N990, N991, N992, N993, N994,
         N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003, N1004,
         N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013, N1014,
         N1015, N1016;
  wire   [12:9] XTEMP;
  wire   [12:0] DIVISION_HEAD;
  wire   [8:0] DIVISION_REMA;
  wire   [12:0] OPER_A;
  wire   [12:0] OPER_B;
  wire   [12:0] SUM_AB;
  wire   [12:0] ZTEMP;
  wire   [3:2] STEP;

  XOR2X1TF \DP_OP_333_124_4748/U28  ( .A(N78), .B(C2_Z_0), .Y(
        DP_OP_333_124_4748_N29) );
  XOR2X1TF \DP_OP_333_124_4748/U27  ( .A(N78), .B(C2_Z_1), .Y(
        DP_OP_333_124_4748_N28) );
  XOR2X1TF \DP_OP_333_124_4748/U26  ( .A(N78), .B(C2_Z_2), .Y(
        DP_OP_333_124_4748_N27) );
  XOR2X1TF \DP_OP_333_124_4748/U25  ( .A(N78), .B(C2_Z_3), .Y(
        DP_OP_333_124_4748_N26) );
  XOR2X1TF \DP_OP_333_124_4748/U24  ( .A(N125), .B(C2_Z_4), .Y(
        DP_OP_333_124_4748_N25) );
  XOR2X1TF \DP_OP_333_124_4748/U23  ( .A(N78), .B(C2_Z_5), .Y(
        DP_OP_333_124_4748_N24) );
  XOR2X1TF \DP_OP_333_124_4748/U22  ( .A(N125), .B(C2_Z_6), .Y(
        DP_OP_333_124_4748_N23) );
  XOR2X1TF \DP_OP_333_124_4748/U21  ( .A(N78), .B(C2_Z_7), .Y(
        DP_OP_333_124_4748_N22) );
  XOR2X1TF \DP_OP_333_124_4748/U20  ( .A(N125), .B(C2_Z_8), .Y(
        DP_OP_333_124_4748_N21) );
  XOR2X1TF \DP_OP_333_124_4748/U19  ( .A(N78), .B(C2_Z_9), .Y(
        DP_OP_333_124_4748_N20) );
  XOR2X1TF \DP_OP_333_124_4748/U18  ( .A(N125), .B(C2_Z_10), .Y(
        DP_OP_333_124_4748_N19) );
  XOR2X1TF \DP_OP_333_124_4748/U17  ( .A(N78), .B(C2_Z_11), .Y(
        DP_OP_333_124_4748_N18) );
  CMPR32X2TF \DP_OP_333_124_4748/U13  ( .A(DP_OP_333_124_4748_N57), .B(N78), 
        .C(DP_OP_333_124_4748_N29), .CO(DP_OP_333_124_4748_N12), .S(
        C152_DATA4_0) );
  ADDHXLTF \DP_OP_333_124_4748/U12  ( .A(DP_OP_333_124_4748_N28), .B(
        DP_OP_333_124_4748_N12), .CO(DP_OP_333_124_4748_N11), .S(C152_DATA4_1)
         );
  ADDHXLTF \DP_OP_333_124_4748/U11  ( .A(DP_OP_333_124_4748_N27), .B(
        DP_OP_333_124_4748_N11), .CO(DP_OP_333_124_4748_N10), .S(C152_DATA4_2)
         );
  ADDHXLTF \DP_OP_333_124_4748/U10  ( .A(DP_OP_333_124_4748_N26), .B(
        DP_OP_333_124_4748_N10), .CO(DP_OP_333_124_4748_N9), .S(C152_DATA4_3)
         );
  ADDHXLTF \DP_OP_333_124_4748/U9  ( .A(DP_OP_333_124_4748_N25), .B(
        DP_OP_333_124_4748_N9), .CO(DP_OP_333_124_4748_N8), .S(C152_DATA4_4)
         );
  ADDHXLTF \DP_OP_333_124_4748/U8  ( .A(DP_OP_333_124_4748_N24), .B(
        DP_OP_333_124_4748_N8), .CO(DP_OP_333_124_4748_N7), .S(C152_DATA4_5)
         );
  ADDHXLTF \DP_OP_333_124_4748/U7  ( .A(DP_OP_333_124_4748_N23), .B(
        DP_OP_333_124_4748_N7), .CO(DP_OP_333_124_4748_N6), .S(C152_DATA4_6)
         );
  ADDHXLTF \DP_OP_333_124_4748/U6  ( .A(DP_OP_333_124_4748_N22), .B(
        DP_OP_333_124_4748_N6), .CO(DP_OP_333_124_4748_N5), .S(C152_DATA4_7)
         );
  ADDHXLTF \DP_OP_333_124_4748/U5  ( .A(DP_OP_333_124_4748_N21), .B(
        DP_OP_333_124_4748_N5), .CO(DP_OP_333_124_4748_N4), .S(C152_DATA4_8)
         );
  ADDHXLTF \DP_OP_333_124_4748/U4  ( .A(DP_OP_333_124_4748_N20), .B(
        DP_OP_333_124_4748_N4), .CO(DP_OP_333_124_4748_N3), .S(C152_DATA4_9)
         );
  ADDHXLTF \DP_OP_333_124_4748/U3  ( .A(DP_OP_333_124_4748_N19), .B(
        DP_OP_333_124_4748_N3), .CO(DP_OP_333_124_4748_N2), .S(C152_DATA4_10)
         );
  ADDHXLTF \DP_OP_333_124_4748/U2  ( .A(DP_OP_333_124_4748_N18), .B(
        DP_OP_333_124_4748_N2), .CO(DP_OP_333_124_4748_N1), .S(C152_DATA4_11)
         );
  CMPR32X2TF \intadd_0/U8  ( .A(X_IN[1]), .B(DIVISION_HEAD[5]), .C(INTADD_0_CI), .CO(INTADD_0_N7), .S(\INTADD_0_SUM[0] ) );
  CMPR32X2TF \intadd_0/U7  ( .A(X_IN[2]), .B(DIVISION_HEAD[6]), .C(INTADD_0_N7), .CO(INTADD_0_N6), .S(\INTADD_0_SUM[1] ) );
  CMPR32X2TF \intadd_0/U6  ( .A(X_IN[3]), .B(DIVISION_HEAD[7]), .C(INTADD_0_N6), .CO(INTADD_0_N5), .S(\INTADD_0_SUM[2] ) );
  CMPR32X2TF \intadd_0/U5  ( .A(X_IN[4]), .B(DIVISION_HEAD[8]), .C(INTADD_0_N5), .CO(INTADD_0_N4), .S(\INTADD_0_SUM[3] ) );
  CMPR32X2TF \intadd_0/U4  ( .A(X_IN[5]), .B(DIVISION_HEAD[9]), .C(INTADD_0_N4), .CO(INTADD_0_N3), .S(\INTADD_0_SUM[4] ) );
  CMPR32X2TF \intadd_0/U3  ( .A(X_IN[6]), .B(DIVISION_HEAD[10]), .C(
        INTADD_0_N3), .CO(INTADD_0_N2), .S(\INTADD_0_SUM[5] ) );
  CMPR32X2TF \intadd_0/U2  ( .A(X_IN[7]), .B(DIVISION_HEAD[11]), .C(
        INTADD_0_N2), .CO(INTADD_0_N1), .S(\INTADD_0_SUM[6] ) );
  DFFSX2TF pre_work_reg ( .D(N695), .CK(CLK), .SN(RST_N), .Q(PRE_WORK), .QN(
        N174) );
  DFFRX2TF \ytemp_reg[10]  ( .D(N684), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[1]), .QN(N172) );
  DFFRX2TF \xtemp_reg[12]  ( .D(N723), .CK(CLK), .RN(RST_N), .Q(XTEMP[12]), 
        .QN(N170) );
  DFFRX2TF \ytemp_reg[9]  ( .D(N685), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[0]), .QN(N167) );
  DFFRX2TF \ytemp_reg[7]  ( .D(N687), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[7]), .QN(N166) );
  DFFRX2TF \ytemp_reg[5]  ( .D(N689), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[5]), .QN(N165) );
  DFFRX2TF \ytemp_reg[3]  ( .D(N691), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[3]), .QN(N164) );
  DFFRX2TF \ytemp_reg[11]  ( .D(N683), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[2]), .QN(N161) );
  DFFRX2TF \xtemp_reg[11]  ( .D(N708), .CK(CLK), .RN(RST_N), .Q(XTEMP[11]), 
        .QN(N154) );
  DFFRX2TF \xtemp_reg[2]  ( .D(N717), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[6]), .QN(N150) );
  DFFRX2TF \ytemp_reg[12]  ( .D(N706), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[3]), .QN(N147) );
  DFFRX2TF \xtemp_reg[10]  ( .D(N709), .CK(CLK), .RN(RST_N), .Q(XTEMP[10]), 
        .QN(N146) );
  DFFRX2TF \ytemp_reg[8]  ( .D(N686), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[8]), .QN(N145) );
  DFFRX2TF \xtemp_reg[5]  ( .D(N714), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[9]), .QN(N144) );
  DFFRX2TF \xtemp_reg[3]  ( .D(N716), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[7]), .QN(N143) );
  DFFRX2TF \xtemp_reg[7]  ( .D(N712), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[11]), .QN(N141) );
  ADDHX1TF \add_x_132_1/U14  ( .A(OPER_B[0]), .B(OPER_A[0]), .CO(
        ADD_X_132_1_N13), .S(SUM_AB[0]) );
  CMPR32X2TF \add_x_132_1/U4  ( .A(OPER_A[10]), .B(OPER_B[10]), .C(
        ADD_X_132_1_N4), .CO(ADD_X_132_1_N3), .S(SUM_AB[10]) );
  CMPR32X2TF \add_x_132_1/U6  ( .A(OPER_A[8]), .B(OPER_B[8]), .C(
        ADD_X_132_1_N6), .CO(ADD_X_132_1_N5), .S(SUM_AB[8]) );
  CMPR32X2TF \add_x_132_1/U10  ( .A(OPER_A[4]), .B(OPER_B[4]), .C(
        ADD_X_132_1_N10), .CO(ADD_X_132_1_N9), .S(SUM_AB[4]) );
  CMPR32X2TF \add_x_132_1/U13  ( .A(OPER_A[1]), .B(OPER_B[1]), .C(
        ADD_X_132_1_N13), .CO(ADD_X_132_1_N12), .S(SUM_AB[1]) );
  CMPR32X2TF \add_x_132_1/U5  ( .A(OPER_A[9]), .B(OPER_B[9]), .C(
        ADD_X_132_1_N5), .CO(ADD_X_132_1_N4), .S(SUM_AB[9]) );
  CMPR32X2TF \add_x_132_1/U12  ( .A(OPER_A[2]), .B(OPER_B[2]), .C(
        ADD_X_132_1_N12), .CO(ADD_X_132_1_N11), .S(SUM_AB[2]) );
  CMPR32X2TF \add_x_132_1/U11  ( .A(OPER_A[3]), .B(OPER_B[3]), .C(
        ADD_X_132_1_N11), .CO(ADD_X_132_1_N10), .S(SUM_AB[3]) );
  CMPR32X2TF \add_x_132_1/U9  ( .A(OPER_A[5]), .B(OPER_B[5]), .C(
        ADD_X_132_1_N9), .CO(ADD_X_132_1_N8), .S(SUM_AB[5]) );
  CMPR32X2TF \add_x_132_1/U3  ( .A(OPER_A[11]), .B(OPER_B[11]), .C(
        ADD_X_132_1_N3), .CO(ADD_X_132_1_N2), .S(SUM_AB[11]) );
  DFFRX1TF \rsht_bits_reg[2]  ( .D(N701), .CK(CLK), .RN(RST_N), .QN(N90) );
  DFFRX1TF \ztemp_reg[0]  ( .D(N669), .CK(CLK), .RN(RST_N), .Q(ZTEMP[0]) );
  DFFRX1TF \wtemp_reg[6]  ( .D(N676), .CK(CLK), .RN(RST_N), .Q(OPER_B[6]) );
  DFFRX1TF \ztemp_reg[6]  ( .D(N663), .CK(CLK), .RN(RST_N), .Q(ZTEMP[6]) );
  DFFRX1TF \ztemp_reg[4]  ( .D(N665), .CK(CLK), .RN(RST_N), .Q(ZTEMP[4]) );
  DFFRX1TF \ztemp_reg[2]  ( .D(N667), .CK(CLK), .RN(RST_N), .Q(ZTEMP[2]) );
  DFFRX1TF \ztemp_reg[1]  ( .D(N668), .CK(CLK), .RN(RST_N), .Q(ZTEMP[1]) );
  DFFRX1TF \ztemp_reg[5]  ( .D(N664), .CK(CLK), .RN(RST_N), .Q(ZTEMP[5]) );
  DFFRX1TF \ztemp_reg[3]  ( .D(N666), .CK(CLK), .RN(RST_N), .Q(ZTEMP[3]) );
  DFFRX1TF \ztemp_reg[7]  ( .D(N662), .CK(CLK), .RN(RST_N), .Q(ZTEMP[7]) );
  DFFRX1TF \ztemp_reg[8]  ( .D(N661), .CK(CLK), .RN(RST_N), .Q(ZTEMP[8]) );
  DFFRX1TF \ztemp_reg[9]  ( .D(N660), .CK(CLK), .RN(RST_N), .Q(ZTEMP[9]) );
  DFFRX1TF \wtemp_reg[5]  ( .D(N677), .CK(CLK), .RN(RST_N), .Q(OPER_B[5]) );
  DFFRX1TF \wtemp_reg[7]  ( .D(N675), .CK(CLK), .RN(RST_N), .Q(OPER_B[7]) );
  DFFRX1TF \ztemp_reg[10]  ( .D(N659), .CK(CLK), .RN(RST_N), .Q(ZTEMP[10]) );
  DFFRX1TF \ztemp_reg[11]  ( .D(N658), .CK(CLK), .RN(RST_N), .Q(ZTEMP[11]) );
  DFFRX1TF \ztemp_reg[12]  ( .D(N657), .CK(CLK), .RN(RST_N), .Q(ZTEMP[12]) );
  DFFRX2TF sign_y_reg ( .D(N694), .CK(CLK), .RN(RST_N), .Q(SIGN_Y), .QN(N177)
         );
  DFFRX2TF \step_reg[2]  ( .D(N696), .CK(CLK), .RN(RST_N), .Q(STEP[2]), .QN(
        N140) );
  DFFRX2TF \step_reg[1]  ( .D(N700), .CK(CLK), .RN(RST_N), .Q(N148), .QN(N121)
         );
  DFFRX2TF \step_reg[3]  ( .D(N721), .CK(CLK), .RN(RST_N), .Q(STEP[3]), .QN(
        N149) );
  DFFRX2TF \step_reg[0]  ( .D(N697), .CK(CLK), .RN(RST_N), .Q(N163), .QN(N122)
         );
  DFFRX2TF SEL_SRC_reg ( .D(N720), .CK(CLK), .RN(RST_N), .Q(POST_WORK), .QN(
        N162) );
  DFFRX2TF \rsht_bits_reg[1]  ( .D(N702), .CK(CLK), .RN(RST_N), .Q(N157), .QN(
        N91) );
  DFFRX2TF \rsht_bits_reg[0]  ( .D(N703), .CK(CLK), .RN(RST_N), .Q(N179), .QN(
        N92) );
  DFFRX2TF SEL_Z_reg ( .D(N670), .CK(CLK), .RN(RST_N), .Q(N169), .QN(N123) );
  DFFRX2TF \rsht_bits_reg[3]  ( .D(N704), .CK(CLK), .RN(RST_N), .Q(
        \RSHT_BITS[3] ), .QN(N188) );
  DFFRX2TF \index_reg[1]  ( .D(N699), .CK(CLK), .RN(RST_N), .Q(N180), .QN(N128) );
  DFFRX2TF \ytemp_reg[0]  ( .D(N705), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[0]), .QN(N178) );
  DFFRX2TF \index_reg[3]  ( .D(N725), .CK(CLK), .RN(RST_N), .Q(N185), .QN(N124) );
  DFFRX2TF \index_reg[0]  ( .D(N726), .CK(CLK), .RN(RST_N), .Q(N156), .QN(N129) );
  DFFRX2TF \wtemp_reg[2]  ( .D(N680), .CK(CLK), .RN(RST_N), .Q(OPER_B[2]), 
        .QN(N155) );
  DFFRX2TF \wtemp_reg[8]  ( .D(N674), .CK(CLK), .RN(RST_N), .Q(OPER_B[8]), 
        .QN(N159) );
  DFFRX2TF \wtemp_reg[0]  ( .D(N682), .CK(CLK), .RN(RST_N), .Q(OPER_B[0]), 
        .QN(N183) );
  DFFRX2TF \wtemp_reg[12]  ( .D(N724), .CK(CLK), .RN(RST_N), .Q(OPER_B[12]), 
        .QN(N186) );
  DFFRX2TF \xtemp_reg[0]  ( .D(N719), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[4]), .QN(N151) );
  DFFRX2TF \wtemp_reg[10]  ( .D(N672), .CK(CLK), .RN(RST_N), .Q(OPER_B[10]), 
        .QN(N160) );
  DFFRX2TF \wtemp_reg[1]  ( .D(N681), .CK(CLK), .RN(RST_N), .Q(OPER_B[1]), 
        .QN(N181) );
  DFFRX2TF \wtemp_reg[4]  ( .D(N678), .CK(CLK), .RN(RST_N), .Q(OPER_B[4]), 
        .QN(N176) );
  DFFRX2TF \wtemp_reg[9]  ( .D(N673), .CK(CLK), .RN(RST_N), .Q(OPER_B[9]), 
        .QN(N187) );
  DFFRX2TF \wtemp_reg[11]  ( .D(N671), .CK(CLK), .RN(RST_N), .Q(OPER_B[11]), 
        .QN(N184) );
  DFFRX2TF \wtemp_reg[3]  ( .D(N679), .CK(CLK), .RN(RST_N), .Q(OPER_B[3]), 
        .QN(N182) );
  DFFRX2TF \ytemp_reg[6]  ( .D(N688), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[6]), .QN(N173) );
  DFFRX2TF \xtemp_reg[4]  ( .D(N715), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[8]), .QN(N152) );
  DFFRX2TF \xtemp_reg[1]  ( .D(N718), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[5]), .QN(N142) );
  DFFRX2TF \xtemp_reg[8]  ( .D(N711), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[12]), .QN(N175) );
  DFFRX2TF \xtemp_reg[6]  ( .D(N713), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[10]), .QN(N153) );
  DFFRX2TF \ytemp_reg[1]  ( .D(N693), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[1]), .QN(N158) );
  DFFRX2TF \ytemp_reg[2]  ( .D(N692), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[2]), .QN(N171) );
  DFFRX2TF \ytemp_reg[4]  ( .D(N690), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[4]), .QN(N168) );
  DFFRX2TF XOR_SRC_reg ( .D(N707), .CK(CLK), .RN(RST_N), .Q(N56), .QN(N73) );
  DFFRX2TF \xtemp_reg[9]  ( .D(N710), .CK(CLK), .RN(RST_N), .Q(XTEMP[9]), .QN(
        N525) );
  DFFRX2TF sign_x_reg ( .D(N722), .CK(CLK), .RN(RST_N), .Q(N962), .QN(N74) );
  DFFRX2TF \index_reg[2]  ( .D(N698), .CK(CLK), .RN(RST_N), .Q(\INDEX[2] ) );
  NAND2X1TF U3 ( .A(ALU_START), .B(N260), .Y(N596) );
  NOR2X1TF U4 ( .A(N929), .B(OPER_A[11]), .Y(N1) );
  XNOR2X1TF U5 ( .A(OPER_A[12]), .B(N1), .Y(N2) );
  AOI22X1TF U6 ( .A0(N2), .A1(N927), .B0(OPER_A[12]), .B1(N849), .Y(N3) );
  OAI21X1TF U7 ( .A0(N967), .A1(N545), .B0(N133), .Y(N4) );
  XNOR2X1TF U8 ( .A(N4), .B(N78), .Y(N5) );
  XNOR2X1TF U9 ( .A(DP_OP_333_124_4748_N1), .B(N5), .Y(N6) );
  NOR2X1TF U10 ( .A(OPER_B[11]), .B(N932), .Y(N7) );
  OAI31X1TF U11 ( .A0(N106), .A1(N7), .A2(OPER_B[12]), .B0(N820), .Y(N8) );
  AOI211X1TF U12 ( .A0(N105), .A1(N6), .B0(N925), .C0(N8), .Y(N9) );
  OAI31X1TF U13 ( .A0(OPER_B[11]), .A1(N932), .A2(N906), .B0(N862), .Y(N10) );
  AOI32X1TF U14 ( .A0(N120), .A1(OPER_B[12]), .A2(N10), .B0(N219), .B1(
        OPER_B[12]), .Y(N11) );
  NAND4BX1TF U15 ( .AN(N816), .B(N3), .C(N9), .D(N11), .Y(N724) );
  AOI32X1TF U16 ( .A0(N107), .A1(N838), .A2(N931), .B0(N183), .B1(N838), .Y(
        N12) );
  AOI211X1TF U17 ( .A0(C152_DATA4_0), .A1(N105), .B0(N879), .C0(N12), .Y(N13)
         );
  OAI21X1TF U18 ( .A0(N849), .A1(N927), .B0(OPER_A[0]), .Y(N14) );
  OAI211X1TF U19 ( .A0(N181), .A1(N882), .B0(N13), .C0(N14), .Y(N682) );
  AND2X1TF U20 ( .A(N190), .B(ZTEMP[10]), .Y(POUT[10]) );
  OAI222X1TF U21 ( .A0(N87), .A1(N170), .B0(N97), .B1(N146), .C0(N81), .C1(
        N147), .Y(FOUT[10]) );
  NOR3X1TF U22 ( .A(N949), .B(N948), .C(N967), .Y(N15) );
  AOI211XLTF U23 ( .A0(N943), .A1(N947), .B0(N966), .C0(N15), .Y(N16) );
  OAI22X1TF U24 ( .A0(N942), .A1(N112), .B0(N941), .B1(N970), .Y(N17) );
  NOR4XLTF U25 ( .A(N946), .B(N944), .C(N945), .D(N17), .Y(N18) );
  MXI2X1TF U26 ( .A(N16), .B(N123), .S0(N18), .Y(N670) );
  AND2X1TF U27 ( .A(N190), .B(ZTEMP[11]), .Y(POUT[11]) );
  NOR2X1TF U28 ( .A(N98), .B(N154), .Y(FOUT[11]) );
  OAI211X1TF U29 ( .A0(N818), .A1(N374), .B0(N608), .C0(N636), .Y(N19) );
  AOI21XLTF U30 ( .A0(N375), .A1(N817), .B0(N19), .Y(N20) );
  NAND3X1TF U31 ( .A(N376), .B(N539), .C(N20), .Y(N21) );
  OAI22X1TF U32 ( .A0(N636), .A1(N759), .B0(N112), .B1(N377), .Y(N22) );
  OAI21X1TF U33 ( .A0(N22), .A1(N742), .B0(N21), .Y(N23) );
  OAI21X1TF U34 ( .A0(N162), .A1(N21), .B0(N23), .Y(N720) );
  OAI21X1TF U35 ( .A0(N881), .A1(N930), .B0(N928), .Y(N24) );
  AO21X1TF U36 ( .A0(N880), .A1(N933), .B0(N878), .Y(N25) );
  AOI22X1TF U37 ( .A0(OPER_A[7]), .A1(N24), .B0(OPER_B[7]), .B1(N25), .Y(N26)
         );
  OAI31X1TF U38 ( .A0(N880), .A1(N106), .A2(OPER_B[7]), .B0(N26), .Y(N27) );
  AOI211X1TF U39 ( .A0(C152_DATA4_7), .A1(N104), .B0(N205), .C0(N27), .Y(N28)
         );
  NAND3BX1TF U40 ( .AN(OPER_A[7]), .B(N881), .C(N927), .Y(N29) );
  OAI211X1TF U41 ( .A0(N882), .A1(N159), .B0(N28), .C0(N29), .Y(N675) );
  AOI22X1TF U42 ( .A0(DIVISION_HEAD[0]), .A1(N1009), .B0(ZTEMP[0]), .B1(N117), 
        .Y(N30) );
  AOI32XLTF U43 ( .A0(N1016), .A1(N30), .A2(N1007), .B0(N973), .B1(N30), .Y(
        N669) );
  NOR3X1TF U44 ( .A(Y_IN[12]), .B(Y_IN[11]), .C(Y_IN[10]), .Y(N31) );
  CLKINVX1TF U45 ( .A(N439), .Y(N32) );
  AOI22X1TF U46 ( .A0(N316), .A1(N32), .B0(N101), .B1(N733), .Y(N33) );
  OAI21X1TF U47 ( .A0(X_IN[4]), .A1(N315), .B0(N85), .Y(N34) );
  OAI22X1TF U48 ( .A0(N101), .A1(N733), .B0(X_IN[6]), .B1(N656), .Y(N35) );
  AOI31X1TF U49 ( .A0(N317), .A1(N33), .A2(N34), .B0(N35), .Y(N36) );
  AOI21X1TF U50 ( .A0(N656), .A1(X_IN[6]), .B0(N36), .Y(N37) );
  OA22X1TF U51 ( .A0(N38), .A1(N37), .B0(N485), .B1(N192), .Y(N39) );
  AO21X1TF U52 ( .A0(N465), .A1(N37), .B0(Y_IN[4]), .Y(N40) );
  AOI22X1TF U53 ( .A0(N485), .A1(N192), .B0(N39), .B1(N40), .Y(N41) );
  AOI2BB2X1TF U54 ( .B0(X_IN[9]), .B1(N41), .A0N(N499), .A1N(N84), .Y(N42) );
  CLKINVX1TF U55 ( .A(N41), .Y(N43) );
  AO21X1TF U56 ( .A0(N497), .A1(N43), .B0(Y_IN[6]), .Y(N44) );
  AOI22X1TF U57 ( .A0(Y_IN[7]), .A1(N499), .B0(N42), .B1(N44), .Y(N45) );
  AOI222XLTF U58 ( .A0(N757), .A1(X_IN[11]), .B0(N757), .B1(N45), .C0(X_IN[11]), .C1(N45), .Y(N46) );
  OAI21X1TF U59 ( .A0(Y_IN[9]), .A1(N303), .B0(N46), .Y(N47) );
  OAI211X1TF U60 ( .A0(X_IN[12]), .A1(N779), .B0(N31), .C0(N47), .Y(N765) );
  CLKINVX1TF U61 ( .A(X_IN[7]), .Y(N38) );
  AND2X1TF U62 ( .A(N190), .B(ZTEMP[12]), .Y(POUT[12]) );
  NOR2X1TF U63 ( .A(N98), .B(N170), .Y(FOUT[12]) );
  CLKINVX1TF U64 ( .A(N859), .Y(N48) );
  OAI31X1TF U65 ( .A0(OPER_B[5]), .A1(N107), .A2(N48), .B0(N893), .Y(N49) );
  AOI21X1TF U66 ( .A0(C152_DATA4_5), .A1(N105), .B0(N49), .Y(N50) );
  NOR2X1TF U67 ( .A(N930), .B(OPER_A[5]), .Y(N51) );
  AOI22X1TF U68 ( .A0(N860), .A1(N51), .B0(OPER_B[6]), .B1(N858), .Y(N52) );
  OAI21X1TF U69 ( .A0(N859), .A1(N107), .B0(N931), .Y(N53) );
  OAI21X1TF U70 ( .A0(N860), .A1(N930), .B0(N928), .Y(N54) );
  AOI22X1TF U71 ( .A0(OPER_B[5]), .A1(N53), .B0(OPER_A[5]), .B1(N54), .Y(N55)
         );
  NAND4X1TF U72 ( .A(N861), .B(N50), .C(N52), .D(N55), .Y(N677) );
  INVX2TF U73 ( .A(N943), .Y(N111) );
  NAND2X2TF U74 ( .A(SIGN_Y), .B(N962), .Y(N968) );
  INVX2TF U75 ( .A(N123), .Y(N58) );
  AOI22X2TF U76 ( .A0(N73), .A1(DIVISION_HEAD[3]), .B0(XTEMP[12]), .B1(N56), 
        .Y(N347) );
  NAND2X1TF U77 ( .A(N769), .B(N761), .Y(N392) );
  NOR3BX2TF U78 ( .AN(ALU_TYPE[2]), .B(ALU_TYPE[0]), .C(ALU_TYPE[1]), .Y(N260)
         );
  OA21XLTF U79 ( .A0(SUM_AB[12]), .A1(N646), .B0(N112), .Y(N135) );
  NAND2X1TF U80 ( .A(N924), .B(N202), .Y(N218) );
  NAND2XLTF U81 ( .A(N795), .B(SUM_AB[8]), .Y(N421) );
  AOI2BB1X1TF U82 ( .A0N(N960), .A1N(N959), .B0(N958), .Y(N1008) );
  CLKINVX1TF U83 ( .A(SUM_AB[4]), .Y(N386) );
  AO21X1TF U84 ( .A0(N772), .A1(N374), .B0(N818), .Y(N506) );
  CLKBUFX2TF U85 ( .A(N189), .Y(DP_OP_333_124_4748_N43) );
  AND2X2TF U86 ( .A(N123), .B(N243), .Y(N258) );
  AND2XLTF U87 ( .A(\INDEX[2] ), .B(N621), .Y(N312) );
  AND2X2TF U88 ( .A(N190), .B(N73), .Y(N241) );
  AND2X2TF U89 ( .A(N110), .B(N190), .Y(N242) );
  CLKINVX1TF U90 ( .A(N192), .Y(N199) );
  CLKINVX1TF U91 ( .A(N834), .Y(N829) );
  CLKINVX1TF U92 ( .A(N617), .Y(N619) );
  CLKINVX1TF U93 ( .A(Y_IN[6]), .Y(N198) );
  CLKBUFX2TF U94 ( .A(N73), .Y(N969) );
  AOI211X1TF U95 ( .A0(X_IN[3]), .A1(N742), .B0(N437), .C0(N436), .Y(N438) );
  AOI211X1TF U96 ( .A0(X_IN[5]), .A1(N742), .B0(N455), .C0(N454), .Y(N456) );
  AOI211X1TF U97 ( .A0(Y_IN[7]), .A1(N742), .B0(N783), .C0(N782), .Y(N784) );
  OA21XLTF U98 ( .A0(SUM_AB[12]), .A1(N391), .B0(N112), .Y(N502) );
  AND2X2TF U99 ( .A(N892), .B(N917), .Y(N933) );
  INVX1TF U100 ( .A(N895), .Y(N877) );
  AOI21X1TF U101 ( .A0(N762), .A1(N307), .B0(N383), .Y(N379) );
  INVX2TF U102 ( .A(N115), .Y(N116) );
  OAI31X1TF U103 ( .A0(N283), .A1(X_IN[11]), .A2(N544), .B0(N282), .Y(N284) );
  AOI22X1TF U104 ( .A0(X_IN[5]), .A1(N441), .B0(N79), .B1(N99), .Y(N443) );
  OAI21XLTF U105 ( .A0(N310), .A1(N625), .B0(N618), .Y(N311) );
  AOI22X1TF U106 ( .A0(X_IN[12]), .A1(N802), .B0(X_IN[11]), .B1(N131), .Y(N433) );
  AOI22X1TF U107 ( .A0(X_IN[2]), .A1(N131), .B0(X_IN[3]), .B1(N802), .Y(N781)
         );
  AOI211X2TF U108 ( .A0(N567), .A1(N943), .B0(N591), .C0(N566), .Y(N593) );
  AOI22X1TF U109 ( .A0(Y_IN[9]), .A1(N797), .B0(X_IN[4]), .B1(N131), .Y(N798)
         );
  AOI21X1TF U110 ( .A0(N639), .A1(N120), .B0(N638), .Y(N642) );
  INVX1TF U111 ( .A(N401), .Y(N402) );
  OAI31X1TF U112 ( .A0(N561), .A1(N562), .A2(N560), .B0(N120), .Y(N578) );
  AOI32XLTF U113 ( .A0(N817), .A1(N943), .A2(N818), .B0(N634), .B1(N120), .Y(
        N640) );
  AOI22X1TF U114 ( .A0(XTEMP[11]), .A1(N126), .B0(N79), .B1(N441), .Y(N355) );
  NAND3XLTF U115 ( .A(N120), .B(N819), .C(N818), .Y(N629) );
  OAI31XLTF U116 ( .A0(N112), .A1(N163), .A2(N628), .B0(N627), .Y(N633) );
  OR2X2TF U117 ( .A(N383), .B(N759), .Y(N796) );
  OAI2BB2XLTF U118 ( .B0(N757), .B1(N799), .A0N(Y_IN[6]), .A1N(N797), .Y(N774)
         );
  NAND4XLTF U119 ( .A(N608), .B(N607), .C(N606), .D(N605), .Y(N609) );
  AOI22X1TF U120 ( .A0(X_IN[2]), .A1(N441), .B0(X_IN[1]), .B1(N797), .Y(N415)
         );
  AOI22X1TF U121 ( .A0(Y_IN[3]), .A1(N797), .B0(DIVISION_REMA[6]), .B1(N114), 
        .Y(N737) );
  AOI22X1TF U122 ( .A0(N192), .A1(N797), .B0(Y_IN[7]), .B1(N786), .Y(N750) );
  AOI22X1TF U123 ( .A0(Y_IN[1]), .A1(N797), .B0(DIVISION_REMA[4]), .B1(N114), 
        .Y(N727) );
  NAND3BXLTF U124 ( .AN(N378), .B(N772), .C(N635), .Y(N367) );
  OAI211XLTF U125 ( .A0(N967), .A1(N366), .B0(N970), .C0(N597), .Y(N368) );
  INVX1TF U126 ( .A(OPER_A[1]), .Y(N827) );
  INVX1TF U127 ( .A(OPER_A[10]), .Y(N910) );
  AOI22X1TF U128 ( .A0(X_IN[2]), .A1(N797), .B0(X_IN[3]), .B1(N441), .Y(N422)
         );
  INVX1TF U129 ( .A(OPER_A[8]), .Y(N885) );
  INVX1TF U130 ( .A(OPER_A[6]), .Y(N869) );
  INVX1TF U131 ( .A(OPER_A[4]), .Y(N857) );
  INVX1TF U132 ( .A(OPER_A[11]), .Y(N926) );
  AOI22X1TF U133 ( .A0(DIVISION_HEAD[2]), .A1(N114), .B0(Y_IN[8]), .B1(N797), 
        .Y(N790) );
  AOI22X1TF U134 ( .A0(DIVISION_REMA[4]), .A1(N103), .B0(ZTEMP[4]), .B1(N169), 
        .Y(N248) );
  AOI22X1TF U135 ( .A0(DIVISION_REMA[7]), .A1(N103), .B0(ZTEMP[7]), .B1(N169), 
        .Y(N251) );
  INVX2TF U136 ( .A(N742), .Y(N95) );
  AOI22X1TF U137 ( .A0(DIVISION_REMA[6]), .A1(N103), .B0(ZTEMP[6]), .B1(N169), 
        .Y(N250) );
  AOI22X1TF U138 ( .A0(DIVISION_HEAD[1]), .A1(N103), .B0(ZTEMP[10]), .B1(N58), 
        .Y(N254) );
  INVX2TF U139 ( .A(DP_OP_333_124_4748_N43), .Y(N78) );
  AOI22X1TF U140 ( .A0(DIVISION_HEAD[3]), .A1(N103), .B0(ZTEMP[12]), .B1(N58), 
        .Y(N257) );
  AOI22X1TF U141 ( .A0(DIVISION_HEAD[2]), .A1(N103), .B0(ZTEMP[11]), .B1(N58), 
        .Y(N255) );
  AOI22X1TF U142 ( .A0(DIVISION_REMA[0]), .A1(N102), .B0(ZTEMP[0]), .B1(N169), 
        .Y(N244) );
  AOI22X1TF U143 ( .A0(DIVISION_REMA[1]), .A1(N102), .B0(ZTEMP[1]), .B1(N169), 
        .Y(N245) );
  INVX2TF U144 ( .A(N731), .Y(N93) );
  AOI22X1TF U145 ( .A0(DIVISION_REMA[5]), .A1(N103), .B0(ZTEMP[5]), .B1(N169), 
        .Y(N249) );
  AOI22X1TF U146 ( .A0(DIVISION_REMA[3]), .A1(N103), .B0(ZTEMP[3]), .B1(N169), 
        .Y(N247) );
  AOI22X1TF U147 ( .A0(DIVISION_REMA[2]), .A1(N102), .B0(ZTEMP[2]), .B1(N169), 
        .Y(N246) );
  AOI22X1TF U148 ( .A0(DIVISION_HEAD[0]), .A1(N103), .B0(ZTEMP[9]), .B1(N58), 
        .Y(N253) );
  AOI22X1TF U149 ( .A0(DIVISION_REMA[8]), .A1(N103), .B0(ZTEMP[8]), .B1(N169), 
        .Y(N252) );
  OAI21XLTF U150 ( .A0(N967), .A1(N315), .B0(N201), .Y(C2_Z_1) );
  OAI21XLTF U151 ( .A0(N967), .A1(N652), .B0(N201), .Y(C2_Z_0) );
  INVX2TF U152 ( .A(N256), .Y(N102) );
  INVX2TF U153 ( .A(N808), .Y(N113) );
  CLKAND2X2TF U154 ( .A(N643), .B(N636), .Y(N542) );
  NAND2BXLTF U155 ( .AN(DP_OP_333_124_4748_N57), .B(N967), .Y(N202) );
  AND2X2TF U156 ( .A(N380), .B(N352), .Y(N731) );
  AND2X2TF U157 ( .A(N352), .B(DP_OP_333_124_4748_N57), .Y(N742) );
  AND2X2TF U158 ( .A(N343), .B(N220), .Y(N943) );
  INVX1TF U159 ( .A(N343), .Y(N952) );
  NAND2XLTF U160 ( .A(N220), .B(N947), .Y(N530) );
  OR3X1TF U161 ( .A(PRE_WORK), .B(N602), .C(N596), .Y(N498) );
  OR2X2TF U162 ( .A(N349), .B(N596), .Y(N808) );
  OR2X2TF U163 ( .A(N169), .B(N243), .Y(N256) );
  CLKAND2X2TF U164 ( .A(ZTEMP[3]), .B(N134), .Y(POUT[3]) );
  CLKAND2X2TF U165 ( .A(ZTEMP[2]), .B(N134), .Y(POUT[2]) );
  CLKAND2X2TF U166 ( .A(ZTEMP[5]), .B(N134), .Y(POUT[5]) );
  CLKAND2X2TF U167 ( .A(ZTEMP[9]), .B(N134), .Y(POUT[9]) );
  CLKAND2X2TF U168 ( .A(ZTEMP[1]), .B(N134), .Y(POUT[1]) );
  CLKAND2X2TF U169 ( .A(ZTEMP[4]), .B(N134), .Y(POUT[4]) );
  CLKAND2X2TF U170 ( .A(ZTEMP[8]), .B(N190), .Y(POUT[8]) );
  INVX2TF U171 ( .A(N969), .Y(N110) );
  INVX2TF U172 ( .A(N193), .Y(N84) );
  INVX2TF U173 ( .A(N195), .Y(N101) );
  CLKAND2X2TF U174 ( .A(ZTEMP[6]), .B(N190), .Y(POUT[6]) );
  CLKAND2X2TF U175 ( .A(ZTEMP[7]), .B(N190), .Y(POUT[7]) );
  CLKAND2X2TF U176 ( .A(ZTEMP[0]), .B(N190), .Y(POUT[0]) );
  NAND2XLTF U177 ( .A(DIVISION_HEAD[4]), .B(N260), .Y(N223) );
  AOI22X1TF U178 ( .A0(X_IN[11]), .A1(N544), .B0(X_IN[12]), .B1(N800), .Y(N278) );
  INVX2TF U179 ( .A(X_IN[3]), .Y(N194) );
  INVX1TF U180 ( .A(X_IN[2]), .Y(N767) );
  INVX2TF U181 ( .A(X_IN[5]), .Y(N195) );
  INVX2TF U182 ( .A(Y_IN[7]), .Y(N193) );
  INVX2TF U183 ( .A(N299), .Y(N79) );
  INVX2TF U184 ( .A(N242), .Y(N80) );
  INVX2TF U185 ( .A(N242), .Y(N81) );
  INVX2TF U186 ( .A(N1016), .Y(N82) );
  INVX2TF U187 ( .A(N1016), .Y(N83) );
  INVX2TF U188 ( .A(N194), .Y(N85) );
  INVX2TF U189 ( .A(N241), .Y(N86) );
  INVX2TF U190 ( .A(N241), .Y(N87) );
  INVX2TF U191 ( .A(N498), .Y(N88) );
  INVX2TF U192 ( .A(N498), .Y(N89) );
  INVX2TF U193 ( .A(N731), .Y(N94) );
  INVX2TF U194 ( .A(N742), .Y(N96) );
  INVX2TF U195 ( .A(N260), .Y(N97) );
  INVX2TF U196 ( .A(N260), .Y(N98) );
  INVX2TF U197 ( .A(N392), .Y(N99) );
  INVX2TF U198 ( .A(N392), .Y(N100) );
  INVX2TF U199 ( .A(N256), .Y(N103) );
  INVX2TF U200 ( .A(N218), .Y(N104) );
  INVX2TF U201 ( .A(N218), .Y(N105) );
  INVX2TF U202 ( .A(N933), .Y(N106) );
  INVX2TF U203 ( .A(N933), .Y(N107) );
  INVX2TF U204 ( .A(N258), .Y(N108) );
  INVX2TF U205 ( .A(N258), .Y(N109) );
  INVX2TF U206 ( .A(N943), .Y(N112) );
  INVX2TF U207 ( .A(N808), .Y(N114) );
  INVX2TF U208 ( .A(N1008), .Y(N115) );
  INVX2TF U209 ( .A(N115), .Y(N117) );
  INVX2TF U210 ( .A(N506), .Y(N118) );
  INVX2TF U211 ( .A(N506), .Y(N119) );
  INVX2TF U212 ( .A(N111), .Y(N120) );
  INVX2TF U213 ( .A(DP_OP_333_124_4748_N43), .Y(N125) );
  INVX2TF U214 ( .A(N93), .Y(N126) );
  AOI222X4TF U215 ( .A0(N484), .A1(N146), .B0(N484), .B1(N499), .C0(N146), 
        .C1(N499), .Y(N494) );
  NOR2X2TF U216 ( .A(N340), .B(N953), .Y(N352) );
  NOR2X2TF U217 ( .A(N349), .B(N967), .Y(N380) );
  NOR3X2TF U218 ( .A(N111), .B(N601), .C(N628), .Y(N614) );
  INVX2TF U219 ( .A(N502), .Y(N127) );
  INVX2TF U220 ( .A(N502), .Y(N130) );
  INVX2TF U221 ( .A(N796), .Y(N131) );
  INVX2TF U222 ( .A(N796), .Y(N132) );
  NAND2X2TF U223 ( .A(N123), .B(N758), .Y(N451) );
  AOI21X2TF U224 ( .A0(N943), .A1(N916), .B0(N219), .Y(N931) );
  AOI211XLTF U225 ( .A0(N827), .A1(N826), .B0(OPER_A[2]), .C0(N911), .Y(N828)
         );
  OAI32XLTF U226 ( .A0(OPER_A[8]), .A1(N886), .A2(N911), .B0(N885), .B1(N884), 
        .Y(N887) );
  OAI32XLTF U227 ( .A0(OPER_A[10]), .A1(N912), .A2(N911), .B0(N910), .B1(N909), 
        .Y(N913) );
  OAI32XLTF U228 ( .A0(OPER_A[6]), .A1(N870), .A2(N911), .B0(N869), .B1(N868), 
        .Y(N871) );
  INVXLTF U229 ( .A(N911), .Y(N908) );
  INVX2TF U230 ( .A(DP_OP_333_124_4748_N57), .Y(N133) );
  CLKBUFX2TF U231 ( .A(N190), .Y(N134) );
  CLKBUFX2TF U232 ( .A(N259), .Y(N190) );
  NOR3XLTF U233 ( .A(N73), .B(N905), .C(N968), .Y(N816) );
  NAND2X2TF U234 ( .A(N966), .B(N924), .Y(N905) );
  AOI21XLTF U235 ( .A0(N819), .A1(N818), .B0(N817), .Y(N830) );
  INVXLTF U236 ( .A(N817), .Y(N377) );
  NOR3BX4TF U237 ( .AN(N382), .B(N379), .C(N126), .Y(N510) );
  AOI222X4TF U238 ( .A0(XTEMP[9]), .A1(X_IN[9]), .B0(XTEMP[9]), .B1(N475), 
        .C0(X_IN[9]), .C1(N475), .Y(N484) );
  AOI222X4TF U239 ( .A0(N175), .A1(N485), .B0(N175), .B1(N461), .C0(N485), 
        .C1(N461), .Y(N475) );
  OAI31XLTF U240 ( .A0(OPER_A[1]), .A1(N911), .A2(OPER_A[0]), .B0(N832), .Y(
        N833) );
  OAI21X2TF U241 ( .A0(N142), .A1(N108), .B0(N245), .Y(OPER_A[1]) );
  NAND2X2TF U242 ( .A(N758), .B(N58), .Y(N555) );
  NOR2X4TF U243 ( .A(N383), .B(N764), .Y(N802) );
  AOI22XLTF U244 ( .A0(DIVISION_HEAD[5]), .A1(N88), .B0(X_IN[7]), .B1(N802), 
        .Y(N385) );
  AOI22XLTF U245 ( .A0(X_IN[10]), .A1(N131), .B0(X_IN[11]), .B1(N802), .Y(N424) );
  NOR4X2TF U246 ( .A(N644), .B(N944), .C(N368), .D(N367), .Y(N638) );
  NOR2X2TF U247 ( .A(N340), .B(N600), .Y(N562) );
  NOR2BX2TF U248 ( .AN(N540), .B(N380), .Y(N625) );
  INVX2TF U249 ( .A(N135), .Y(N136) );
  INVX2TF U250 ( .A(N135), .Y(N137) );
  AOI22X2TF U251 ( .A0(N347), .A1(N345), .B0(N942), .B1(N348), .Y(N917) );
  CLKBUFX2TF U252 ( .A(N1009), .Y(N138) );
  NOR2X1TF U253 ( .A(N116), .B(N189), .Y(N1009) );
  XNOR2X1TF U254 ( .A(OPER_A[12]), .B(ADD_X_132_1_N2), .Y(N139) );
  CMPR32X2TF U255 ( .A(OPER_A[7]), .B(OPER_B[7]), .C(ADD_X_132_1_N7), .CO(
        ADD_X_132_1_N6), .S(SUM_AB[7]) );
  CMPR32X2TF U256 ( .A(OPER_A[6]), .B(OPER_B[6]), .C(ADD_X_132_1_N8), .CO(
        ADD_X_132_1_N7), .S(SUM_AB[6]) );
  XNOR2X2TF U257 ( .A(N139), .B(OPER_B[12]), .Y(SUM_AB[12]) );
  AOI222XLTF U258 ( .A0(DIVISION_HEAD[1]), .A1(DIVISION_HEAD[0]), .B0(
        DIVISION_HEAD[1]), .B1(N316), .C0(DIVISION_HEAD[0]), .C1(N315), .Y(
        N318) );
  AOI32X1TF U259 ( .A0(N120), .A1(N56), .A2(N560), .B0(N614), .B1(N73), .Y(
        N541) );
  AOI22X1TF U260 ( .A0(N73), .A1(N162), .B0(POST_WORK), .B1(N110), .Y(N243) );
  NAND2X1TF U261 ( .A(N315), .B(N652), .Y(N317) );
  NAND2X1TF U262 ( .A(N474), .B(N473), .Y(N483) );
  NOR2X1TF U263 ( .A(SUM_AB[8]), .B(N459), .Y(N474) );
  NOR2X1TF U264 ( .A(SUM_AB[10]), .B(N483), .Y(N496) );
  OA22X1TF U265 ( .A0(N764), .A1(N554), .B0(N759), .B1(N760), .Y(N307) );
  INVX2TF U266 ( .A(N924), .Y(N219) );
  OAI21X1TF U267 ( .A0(N948), .A1(N606), .B0(N643), .Y(N958) );
  NAND2X1TF U268 ( .A(Y_IN[1]), .B(Y_IN[0]), .Y(N316) );
  NAND2X1TF U269 ( .A(N561), .B(N348), .Y(N911) );
  NOR2X2TF U270 ( .A(N219), .B(N111), .Y(N892) );
  OR2X2TF U271 ( .A(N958), .B(N197), .Y(N924) );
  NOR2X1TF U272 ( .A(\INDEX[2] ), .B(N617), .Y(N310) );
  NAND2X1TF U273 ( .A(N129), .B(N128), .Y(N617) );
  OAI21X1TF U274 ( .A0(DIVISION_HEAD[12]), .A1(N545), .B0(N339), .Y(N948) );
  AOI2BB1X1TF U275 ( .A0N(DIVISION_HEAD[6]), .A1N(N328), .B0(Y_IN[6]), .Y(N326) );
  AOI2BB1X1TF U276 ( .A0N(DIVISION_HEAD[4]), .A1N(N324), .B0(Y_IN[4]), .Y(N322) );
  NAND2X1TF U277 ( .A(PRE_WORK), .B(N125), .Y(N383) );
  AOI211X1TF U278 ( .A0(Y_IN[11]), .A1(N303), .B0(Y_IN[12]), .C0(N284), .Y(
        N762) );
  CLKBUFX2TF U279 ( .A(N967), .Y(N189) );
  NAND2X1TF U280 ( .A(N907), .B(N892), .Y(N928) );
  AOI2BB1X1TF U281 ( .A0N(N604), .A1N(N344), .B0(N959), .Y(N197) );
  NOR2X1TF U282 ( .A(PRE_WORK), .B(N341), .Y(N343) );
  NAND2X1TF U283 ( .A(N122), .B(N148), .Y(N601) );
  NOR2X1TF U284 ( .A(N124), .B(N624), .Y(N341) );
  CLKBUFX2TF U285 ( .A(Y_IN[5]), .Y(N192) );
  NAND2X1TF U286 ( .A(N140), .B(N149), .Y(N340) );
  NAND2X1TF U287 ( .A(N451), .B(N457), .Y(N468) );
  NAND2X2TF U288 ( .A(N543), .B(N382), .Y(N457) );
  CLKBUFX2TF U289 ( .A(N777), .Y(N191) );
  NAND2X1TF U290 ( .A(N121), .B(N122), .Y(N953) );
  AND2X2TF U291 ( .A(ALU_START), .B(N134), .Y(N220) );
  NAND2X1TF U292 ( .A(N562), .B(N380), .Y(N606) );
  NAND2X2TF U293 ( .A(N221), .B(ALU_START), .Y(N967) );
  NAND2X1TF U294 ( .A(N174), .B(N366), .Y(N349) );
  NAND2X1TF U295 ( .A(N124), .B(N310), .Y(N366) );
  NAND2X1TF U296 ( .A(N121), .B(N163), .Y(N600) );
  AND2X2TF U297 ( .A(N196), .B(ALU_TYPE[1]), .Y(N221) );
  AOI211X1TF U298 ( .A0(N220), .A1(N604), .B0(N946), .C0(N603), .Y(N607) );
  NOR3X1TF U299 ( .A(N602), .B(N601), .C(N772), .Y(N603) );
  OR3X1TF U300 ( .A(N876), .B(N875), .C(N214), .Y(N676) );
  OAI2BB2XLTF U301 ( .B0(N877), .B1(N968), .A0N(C152_DATA4_6), .A1N(N105), .Y(
        N214) );
  OAI2BB2XLTF U302 ( .B0(N874), .B1(N919), .A0N(N219), .A1N(OPER_B[6]), .Y(
        N875) );
  INVX2TF U303 ( .A(N457), .Y(N472) );
  AOI32X1TF U304 ( .A0(N966), .A1(N115), .A2(N965), .B0(N120), .B1(N115), .Y(
        N1016) );
  NOR2BX2TF U305 ( .AN(N543), .B(N553), .Y(N809) );
  NOR2X1TF U306 ( .A(N174), .B(N596), .Y(N354) );
  NAND2X1TF U307 ( .A(N957), .B(DP_OP_333_124_4748_N57), .Y(N646) );
  INVX2TF U308 ( .A(N365), .Y(N758) );
  NAND2X1TF U309 ( .A(N380), .B(N957), .Y(N365) );
  NAND2X1TF U310 ( .A(N892), .B(N865), .Y(N882) );
  NOR2X1TF U311 ( .A(N56), .B(N905), .Y(N895) );
  AND2X2TF U312 ( .A(N220), .B(PRE_WORK), .Y(DP_OP_333_124_4748_N57) );
  AOI21X1TF U313 ( .A0(N949), .A1(N964), .B0(N364), .Y(N966) );
  NAND2X1TF U314 ( .A(N140), .B(STEP[3]), .Y(N628) );
  NOR2X2TF U315 ( .A(N340), .B(N601), .Y(N957) );
  NAND2X1TF U316 ( .A(N341), .B(N174), .Y(N346) );
  NAND3X1TF U317 ( .A(N959), .B(N967), .C(N596), .Y(N643) );
  INVX2TF U318 ( .A(N220), .Y(N959) );
  NOR3BX1TF U319 ( .AN(ALU_TYPE[0]), .B(ALU_TYPE[1]), .C(ALU_TYPE[2]), .Y(N259) );
  AO22X1TF U320 ( .A0(N373), .A1(XTEMP[12]), .B0(N361), .B1(N962), .Y(N722) );
  AOI32X1TF U321 ( .A0(N964), .A1(N362), .A2(N955), .B0(N970), .B1(N362), .Y(
        N363) );
  NAND2X1TF U322 ( .A(N947), .B(DP_OP_333_124_4748_N57), .Y(N631) );
  NAND2X1TF U323 ( .A(N639), .B(N114), .Y(N611) );
  NAND2X1TF U324 ( .A(N105), .B(C152_DATA4_8), .Y(N215) );
  AOI32X1TF U325 ( .A0(N118), .A1(DIVISION_HEAD[4]), .A2(N745), .B0(N468), 
        .B1(DIVISION_HEAD[4]), .Y(N389) );
  OAI22X1TF U326 ( .A0(N525), .A1(N94), .B0(N485), .B1(N96), .Y(N486) );
  INVX2TF U327 ( .A(N1012), .Y(N1007) );
  OAI2BB2XLTF U328 ( .B0(N56), .B1(N968), .A0N(N968), .A1N(N56), .Y(N971) );
  NAND2X1TF U329 ( .A(N643), .B(N95), .Y(N945) );
  NAND2X1TF U330 ( .A(N562), .B(DP_OP_333_124_4748_N57), .Y(N391) );
  INVX2TF U331 ( .A(N113), .Y(N772) );
  NOR2X2TF U332 ( .A(N758), .B(N191), .Y(N756) );
  NAND2X1TF U333 ( .A(N352), .B(N113), .Y(N540) );
  NOR2X1TF U334 ( .A(N953), .B(N628), .Y(N560) );
  OAI21X2TF U335 ( .A0(N151), .A1(N108), .B0(N244), .Y(OPER_A[0]) );
  NOR2X1TF U336 ( .A(N601), .B(N951), .Y(N561) );
  NAND2X1TF U337 ( .A(STEP[2]), .B(N149), .Y(N951) );
  OAI32X1TF U338 ( .A0(N645), .A1(N177), .A2(N945), .B0(N147), .B1(N646), .Y(
        N694) );
  OAI21X1TF U339 ( .A0(N174), .A1(N644), .B0(N643), .Y(N695) );
  AOI22X1TF U340 ( .A0(N539), .A1(N73), .B0(N538), .B1(N537), .Y(N707) );
  INVX2TF U341 ( .A(N539), .Y(N537) );
  OAI31X1TF U342 ( .A0(N536), .A1(N535), .A2(N534), .B0(N533), .Y(N538) );
  AOI211X1TF U343 ( .A0(N532), .A1(XTEMP[12]), .B0(N531), .C0(N530), .Y(N533)
         );
  OAI31X1TF U344 ( .A0(DIVISION_HEAD[1]), .A1(N529), .A2(N146), .B0(N528), .Y(
        N532) );
  AOI22X1TF U345 ( .A0(N527), .A1(N526), .B0(XTEMP[11]), .B1(N161), .Y(N528)
         );
  OAI22X1TF U346 ( .A0(DIVISION_HEAD[0]), .A1(N525), .B0(DIVISION_REMA[8]), 
        .B1(N175), .Y(N526) );
  INVX2TF U347 ( .A(N535), .Y(N527) );
  NOR2X1TF U348 ( .A(XTEMP[11]), .B(N161), .Y(N529) );
  OAI22X1TF U349 ( .A0(DIVISION_HEAD[12]), .A1(N145), .B0(XTEMP[12]), .B1(N147), .Y(N534) );
  OAI21X1TF U350 ( .A0(XTEMP[11]), .A1(N161), .B0(N524), .Y(N535) );
  AOI22X1TF U351 ( .A0(DIVISION_HEAD[0]), .A1(N525), .B0(DIVISION_HEAD[1]), 
        .B1(N146), .Y(N524) );
  AOI21X1TF U352 ( .A0(DIVISION_HEAD[11]), .A1(N166), .B0(N523), .Y(N536) );
  AOI211X1TF U353 ( .A0(DIVISION_REMA[6]), .A1(N153), .B0(N522), .C0(N521), 
        .Y(N523) );
  NOR2X1TF U354 ( .A(DIVISION_HEAD[11]), .B(N166), .Y(N521) );
  AOI21X1TF U355 ( .A0(DIVISION_HEAD[9]), .A1(N165), .B0(N519), .Y(N520) );
  AOI211X1TF U356 ( .A0(DIVISION_REMA[4]), .A1(N152), .B0(N518), .C0(N517), 
        .Y(N519) );
  NOR2X1TF U357 ( .A(DIVISION_HEAD[9]), .B(N165), .Y(N517) );
  AOI21X1TF U358 ( .A0(DIVISION_HEAD[7]), .A1(N164), .B0(N515), .Y(N516) );
  AOI211X1TF U359 ( .A0(N514), .A1(DIVISION_REMA[2]), .B0(N513), .C0(N512), 
        .Y(N515) );
  NOR2X1TF U360 ( .A(DIVISION_HEAD[7]), .B(N164), .Y(N513) );
  OAI21X1TF U361 ( .A0(DIVISION_HEAD[5]), .A1(N158), .B0(N511), .Y(N514) );
  OAI211X1TF U362 ( .A0(DIVISION_REMA[1]), .A1(N142), .B0(DIVISION_REMA[0]), 
        .C0(N151), .Y(N511) );
  OAI21X1TF U363 ( .A0(N593), .A1(N582), .B0(N581), .Y(N702) );
  AOI31X1TF U364 ( .A0(N580), .A1(N585), .A2(N587), .B0(N579), .Y(N582) );
  OAI22X1TF U365 ( .A0(N128), .A1(N578), .B0(N589), .B1(N585), .Y(N579) );
  OAI21X1TF U366 ( .A0(N128), .A1(N616), .B0(N615), .Y(N699) );
  AOI31X1TF U367 ( .A0(N614), .A1(N617), .A2(N613), .B0(N612), .Y(N615) );
  OAI32X1TF U368 ( .A0(N625), .A1(N626), .A2(N617), .B0(N613), .B1(N625), .Y(
        N612) );
  AOI22X1TF U369 ( .A0(N593), .A1(N92), .B0(N577), .B1(N576), .Y(N703) );
  AOI211X1TF U370 ( .A0(N591), .A1(N156), .B0(N575), .C0(N786), .Y(N577) );
  AOI21X1TF U371 ( .A0(N574), .A1(N772), .B0(N179), .Y(N575) );
  OAI21X1TF U372 ( .A0(N129), .A1(N616), .B0(N309), .Y(N726) );
  OAI21X1TF U373 ( .A0(N308), .A1(N379), .B0(N616), .Y(N309) );
  AOI32X1TF U374 ( .A0(N625), .A1(N631), .A2(N376), .B0(N156), .B1(N631), .Y(
        N308) );
  OAI31X1TF U375 ( .A0(N626), .A1(N625), .A2(N624), .B0(N623), .Y(N698) );
  AOI22X1TF U376 ( .A0(\INDEX[2] ), .A1(N622), .B0(N621), .B1(N620), .Y(N623)
         );
  OAI21X1TF U377 ( .A0(N619), .A1(N625), .B0(N618), .Y(N622) );
  AOI32X1TF U378 ( .A0(N312), .A1(N124), .A2(N614), .B0(N185), .B1(N311), .Y(
        N314) );
  NOR2X1TF U379 ( .A(N626), .B(N620), .Y(N618) );
  AOI21X1TF U380 ( .A0(\INDEX[2] ), .A1(N621), .B0(N376), .Y(N620) );
  INVX2TF U381 ( .A(N616), .Y(N626) );
  INVX2TF U382 ( .A(N613), .Y(N621) );
  OAI211X1TF U383 ( .A0(N112), .A1(N370), .B0(N641), .C0(N369), .Y(N721) );
  AOI22X1TF U384 ( .A0(STEP[3]), .A1(N638), .B0(N375), .B1(N570), .Y(N369) );
  OAI211X1TF U385 ( .A0(N178), .A1(N611), .B0(N627), .C0(N610), .Y(N700) );
  AOI21X1TF U386 ( .A0(N638), .A1(N148), .B0(N609), .Y(N610) );
  NOR3X1TF U387 ( .A(STEP[3]), .B(N112), .C(N600), .Y(N946) );
  AOI211X1TF U388 ( .A0(N819), .A1(N375), .B0(N373), .C0(N372), .Y(N608) );
  AOI21X1TF U389 ( .A0(N381), .A1(N371), .B0(N772), .Y(N372) );
  NOR2X1TF U390 ( .A(N111), .B(N818), .Y(N375) );
  OAI22X1TF U391 ( .A0(N90), .A1(N594), .B0(N593), .B1(N592), .Y(N701) );
  AOI21X1TF U392 ( .A0(\INDEX[2] ), .A1(N591), .B0(N590), .Y(N592) );
  OAI22X1TF U393 ( .A0(N589), .A1(N588), .B0(N587), .B1(N586), .Y(N590) );
  INVX2TF U394 ( .A(N584), .Y(N589) );
  AOI21X1TF U395 ( .A0(N585), .A1(N584), .B0(N583), .Y(N594) );
  OAI211X1TF U396 ( .A0(N642), .A1(N140), .B0(N641), .C0(N640), .Y(N696) );
  NOR2X1TF U397 ( .A(N645), .B(N363), .Y(N641) );
  OAI21X1TF U398 ( .A0(N352), .A1(N261), .B0(N120), .Y(N362) );
  INVX2TF U399 ( .A(N646), .Y(N645) );
  OAI22X1TF U400 ( .A0(N163), .A1(N951), .B0(N818), .B1(N964), .Y(N634) );
  AOI211X1TF U401 ( .A0(N638), .A1(N163), .B0(N633), .C0(N632), .Y(N637) );
  INVX2TF U402 ( .A(N262), .Y(N630) );
  AOI31X1TF U403 ( .A0(N953), .A1(N371), .A2(N381), .B0(N772), .Y(N262) );
  AOI21X1TF U404 ( .A0(N125), .A1(N599), .B0(N598), .Y(N627) );
  OAI21X1TF U405 ( .A0(N597), .A1(N596), .B0(N595), .Y(N598) );
  OAI22X1TF U406 ( .A0(N593), .A1(N573), .B0(N572), .B1(N188), .Y(N704) );
  AOI21X1TF U407 ( .A0(N588), .A1(N584), .B0(N583), .Y(N572) );
  OAI21X1TF U408 ( .A0(N90), .A1(N587), .B0(N580), .Y(N586) );
  INVX2TF U409 ( .A(N611), .Y(N580) );
  INVX2TF U410 ( .A(N593), .Y(N576) );
  OAI31X1TF U411 ( .A0(N602), .A1(N601), .A2(N772), .B0(N574), .Y(N584) );
  OAI32X1TF U412 ( .A0(N571), .A1(N819), .A2(N570), .B0(N120), .B1(N571), .Y(
        N574) );
  INVX2TF U413 ( .A(N569), .Y(N571) );
  AOI21X1TF U414 ( .A0(N591), .A1(N185), .B0(N568), .Y(N573) );
  AOI32X1TF U415 ( .A0(N562), .A1(N114), .A2(N178), .B0(N957), .B1(N113), .Y(
        N564) );
  AOI31X1TF U416 ( .A0(N120), .A1(N819), .A2(N818), .B0(N945), .Y(N565) );
  INVX2TF U417 ( .A(N578), .Y(N591) );
  AOI22X1TF U418 ( .A0(N891), .A1(N892), .B0(N219), .B1(OPER_B[8]), .Y(N216)
         );
  OAI21X1TF U419 ( .A0(N890), .A1(N159), .B0(N889), .Y(N891) );
  AOI211X1TF U420 ( .A0(N915), .A1(OPER_B[9]), .B0(N888), .C0(N887), .Y(N889)
         );
  AOI21X1TF U421 ( .A0(N908), .A1(N886), .B0(N907), .Y(N884) );
  NOR3X1TF U422 ( .A(N906), .B(OPER_B[8]), .C(N883), .Y(N888) );
  AOI21X1TF U423 ( .A0(N883), .A1(N917), .B0(N916), .Y(N890) );
  OAI211X1TF U424 ( .A0(N1007), .A1(N982), .B0(N981), .C0(N980), .Y(N666) );
  AOI22X1TF U425 ( .A0(DIVISION_HEAD[3]), .A1(N138), .B0(ZTEMP[3]), .B1(N117), 
        .Y(N981) );
  OAI211X1TF U426 ( .A0(N1007), .A1(N994), .B0(N993), .C0(N992), .Y(N662) );
  AOI22X1TF U427 ( .A0(DIVISION_HEAD[7]), .A1(N1009), .B0(ZTEMP[7]), .B1(N117), 
        .Y(N993) );
  OAI211X1TF U428 ( .A0(N1007), .A1(N988), .B0(N987), .C0(N986), .Y(N664) );
  AOI22X1TF U429 ( .A0(DIVISION_HEAD[5]), .A1(N138), .B0(ZTEMP[5]), .B1(N117), 
        .Y(N987) );
  AOI22X1TF U430 ( .A0(SUM_AB[1]), .A1(N82), .B0(N974), .B1(N1012), .Y(N975)
         );
  AOI22X1TF U431 ( .A0(DIVISION_HEAD[1]), .A1(N138), .B0(ZTEMP[1]), .B1(N116), 
        .Y(N976) );
  AOI22X1TF U432 ( .A0(SUM_AB[2]), .A1(N82), .B0(N977), .B1(N1012), .Y(N978)
         );
  AOI22X1TF U433 ( .A0(DIVISION_HEAD[2]), .A1(N138), .B0(ZTEMP[2]), .B1(N116), 
        .Y(N979) );
  AOI22X1TF U434 ( .A0(SUM_AB[4]), .A1(N82), .B0(N983), .B1(N1012), .Y(N984)
         );
  AOI22X1TF U435 ( .A0(DIVISION_HEAD[4]), .A1(N138), .B0(ZTEMP[4]), .B1(N117), 
        .Y(N985) );
  AOI22X1TF U436 ( .A0(SUM_AB[6]), .A1(N82), .B0(N989), .B1(N1012), .Y(N990)
         );
  AOI22X1TF U437 ( .A0(DIVISION_HEAD[6]), .A1(N138), .B0(ZTEMP[6]), .B1(N117), 
        .Y(N991) );
  OAI21X1TF U438 ( .A0(N447), .A1(N446), .B0(N457), .Y(N448) );
  AOI22X1TF U439 ( .A0(DIVISION_HEAD[11]), .A1(N89), .B0(X_IN[12]), .B1(N132), 
        .Y(N442) );
  AOI22X1TF U440 ( .A0(SUM_AB[6]), .A1(N127), .B0(N490), .B1(N989), .Y(N444)
         );
  OAI22X1TF U441 ( .A0(N144), .A1(N94), .B0(N439), .B1(N96), .Y(N447) );
  AOI22X1TF U442 ( .A0(SUM_AB[8]), .A1(N82), .B0(N995), .B1(N1012), .Y(N996)
         );
  AOI22X1TF U443 ( .A0(DIVISION_HEAD[8]), .A1(N138), .B0(ZTEMP[8]), .B1(N116), 
        .Y(N997) );
  OAI211X1TF U444 ( .A0(N1007), .A1(N1000), .B0(N999), .C0(N998), .Y(N660) );
  AOI22X1TF U445 ( .A0(DIVISION_HEAD[9]), .A1(N1009), .B0(ZTEMP[9]), .B1(N117), 
        .Y(N999) );
  INVX2TF U446 ( .A(N876), .Y(N213) );
  AOI31X1TF U447 ( .A0(N837), .A1(N836), .A2(N835), .B0(N919), .Y(N839) );
  AOI32X1TF U448 ( .A0(N834), .A1(OPER_B[2]), .A2(N917), .B0(N916), .B1(
        OPER_B[2]), .Y(N835) );
  AOI22X1TF U449 ( .A0(N915), .A1(OPER_B[3]), .B0(OPER_A[2]), .B1(N833), .Y(
        N836) );
  AOI31X1TF U450 ( .A0(N917), .A1(N155), .A2(N829), .B0(N828), .Y(N837) );
  AOI211X1TF U451 ( .A0(N219), .A1(OPER_B[10]), .B0(N922), .C0(N923), .Y(N217)
         );
  AOI21X1TF U452 ( .A0(N972), .A1(N968), .B0(N905), .Y(N923) );
  AOI21X1TF U453 ( .A0(N921), .A1(N920), .B0(N919), .Y(N922) );
  AOI32X1TF U454 ( .A0(N918), .A1(OPER_B[10]), .A2(N917), .B0(N916), .B1(
        OPER_B[10]), .Y(N920) );
  AOI211X1TF U455 ( .A0(N915), .A1(OPER_B[11]), .B0(N914), .C0(N913), .Y(N921)
         );
  AOI21X1TF U456 ( .A0(N908), .A1(N912), .B0(N907), .Y(N909) );
  NOR3X1TF U457 ( .A(N906), .B(OPER_B[10]), .C(N918), .Y(N914) );
  OAI22X1TF U458 ( .A0(N472), .A1(N471), .B0(N470), .B1(N175), .Y(N711) );
  AOI211X1TF U459 ( .A0(N995), .A1(N490), .B0(N467), .C0(N466), .Y(N471) );
  OAI211X1TF U460 ( .A0(N465), .A1(N605), .B0(N464), .C0(N463), .Y(N466) );
  AOI22X1TF U461 ( .A0(XTEMP[9]), .A1(N89), .B0(N795), .B1(SUM_AB[12]), .Y(
        N463) );
  NOR2X1TF U462 ( .A(DIVISION_HEAD[12]), .B(N469), .Y(N462) );
  AOI22X1TF U463 ( .A0(X_IN[8]), .A1(N461), .B0(INTADD_0_N1), .B1(N485), .Y(
        N469) );
  OAI22X1TF U464 ( .A0(N141), .A1(N94), .B0(N460), .B1(N96), .Y(N467) );
  AOI211X1TF U465 ( .A0(OPER_B[6]), .A1(N873), .B0(N872), .C0(N871), .Y(N874)
         );
  AOI21X1TF U466 ( .A0(N908), .A1(N870), .B0(N907), .Y(N868) );
  OAI31X1TF U467 ( .A0(N906), .A1(OPER_B[6]), .A2(N867), .B0(N866), .Y(N872)
         );
  AOI21X1TF U468 ( .A0(OPER_B[7]), .A1(N865), .B0(N864), .Y(N866) );
  OAI21X1TF U469 ( .A0(N906), .A1(N863), .B0(N862), .Y(N873) );
  AOI32X1TF U470 ( .A0(N390), .A1(N389), .A2(N388), .B0(N472), .B1(N389), .Y(
        N719) );
  OAI211X1TF U471 ( .A0(N386), .A1(N555), .B0(N385), .C0(N384), .Y(N387) );
  AOI22X1TF U472 ( .A0(X_IN[6]), .A1(N132), .B0(X_IN[5]), .B1(N100), .Y(N384)
         );
  AOI22X1TF U473 ( .A0(DIVISION_HEAD[3]), .A1(N731), .B0(SUM_AB[0]), .B1(N378), 
        .Y(N390) );
  AOI32X1TF U474 ( .A0(N409), .A1(N457), .A2(N408), .B0(N472), .B1(N150), .Y(
        N717) );
  AOI211X1TF U475 ( .A0(DIVISION_HEAD[7]), .A1(N89), .B0(N407), .C0(N406), .Y(
        N408) );
  OAI211X1TF U476 ( .A0(N96), .A1(N745), .B0(N405), .C0(N404), .Y(N406) );
  AOI21X1TF U477 ( .A0(N490), .A1(N977), .B0(N403), .Y(N404) );
  OAI22X1TF U478 ( .A0(N142), .A1(N93), .B0(N150), .B1(N451), .Y(N403) );
  AOI22X1TF U479 ( .A0(X_IN[1]), .A1(N441), .B0(N795), .B1(SUM_AB[6]), .Y(N405) );
  OAI21X1TF U480 ( .A0(N497), .A1(N744), .B0(N400), .Y(N407) );
  AOI22X1TF U481 ( .A0(X_IN[8]), .A1(N132), .B0(X_IN[7]), .B1(N100), .Y(N400)
         );
  AOI32X1TF U482 ( .A0(N428), .A1(N457), .A2(N427), .B0(N472), .B1(N152), .Y(
        N715) );
  AOI211X1TF U483 ( .A0(N490), .A1(N983), .B0(N426), .C0(N425), .Y(N427) );
  AOI22X1TF U484 ( .A0(DIVISION_HEAD[9]), .A1(N88), .B0(X_IN[9]), .B1(N100), 
        .Y(N423) );
  OAI22X1TF U485 ( .A0(N143), .A1(N94), .B0(N152), .B1(N451), .Y(N426) );
  AOI32X1TF U486 ( .A0(N399), .A1(N457), .A2(N398), .B0(N472), .B1(N142), .Y(
        N718) );
  AOI211X1TF U487 ( .A0(N490), .A1(N974), .B0(N397), .C0(N396), .Y(N398) );
  OAI211X1TF U488 ( .A0(N555), .A1(N429), .B0(N395), .C0(N394), .Y(N396) );
  AOI21X1TF U489 ( .A0(DIVISION_HEAD[4]), .A1(N731), .B0(N393), .Y(N394) );
  OAI22X1TF U490 ( .A0(N142), .A1(N451), .B0(N745), .B1(N605), .Y(N393) );
  AOI22X1TF U491 ( .A0(DIVISION_HEAD[6]), .A1(N89), .B0(X_IN[7]), .B1(N131), 
        .Y(N395) );
  OAI22X1TF U492 ( .A0(N460), .A1(N392), .B0(N485), .B1(N744), .Y(N397) );
  OAI22X1TF U493 ( .A0(N510), .A1(N482), .B0(N481), .B1(N525), .Y(N710) );
  AOI211X1TF U494 ( .A0(SUM_AB[9]), .A1(N130), .B0(N479), .C0(N478), .Y(N482)
         );
  OAI211X1TF U495 ( .A0(N1000), .A1(N504), .B0(N477), .C0(N476), .Y(N478) );
  AOI22X1TF U496 ( .A0(XTEMP[10]), .A1(N89), .B0(X_IN[7]), .B1(N797), .Y(N477)
         );
  OAI22X1TF U497 ( .A0(N175), .A1(N94), .B0(N485), .B1(N605), .Y(N479) );
  AOI32X1TF U498 ( .A0(N458), .A1(N457), .A2(N456), .B0(N472), .B1(N141), .Y(
        N712) );
  OAI211X1TF U499 ( .A0(N504), .A1(N994), .B0(N453), .C0(N452), .Y(N454) );
  AOI22X1TF U500 ( .A0(DIVISION_HEAD[12]), .A1(N88), .B0(X_IN[12]), .B1(N99), 
        .Y(N452) );
  AOI22X1TF U501 ( .A0(DIVISION_HEAD[11]), .A1(N801), .B0(DIVISION_HEAD[10]), 
        .B1(N126), .Y(N453) );
  OAI22X1TF U502 ( .A0(N460), .A1(N605), .B0(N555), .B1(N495), .Y(N455) );
  AOI22X1TF U503 ( .A0(SUM_AB[10]), .A1(N83), .B0(N1001), .B1(N1012), .Y(N1002) );
  AOI22X1TF U504 ( .A0(DIVISION_HEAD[10]), .A1(N138), .B0(ZTEMP[10]), .B1(N117), .Y(N1003) );
  AOI32X1TF U505 ( .A0(N794), .A1(N811), .A2(N793), .B0(N809), .B1(N172), .Y(
        N684) );
  AOI21X1TF U506 ( .A0(N792), .A1(N1001), .B0(N791), .Y(N793) );
  AOI22X1TF U507 ( .A0(X_IN[2]), .A1(N100), .B0(X_IN[4]), .B1(N802), .Y(N787)
         );
  AOI22X1TF U508 ( .A0(DIVISION_HEAD[0]), .A1(N126), .B0(DIVISION_HEAD[1]), 
        .B1(N801), .Y(N788) );
  AOI22X1TF U509 ( .A0(Y_IN[10]), .A1(N786), .B0(X_IN[3]), .B1(N132), .Y(N789)
         );
  AOI22X1TF U510 ( .A0(N795), .A1(SUM_AB[1]), .B0(SUM_AB[10]), .B1(N137), .Y(
        N794) );
  OAI22X1TF U511 ( .A0(N510), .A1(N493), .B0(N492), .B1(N146), .Y(N709) );
  AOI21X1TF U512 ( .A0(N490), .A1(N1001), .B0(N489), .Y(N493) );
  OAI211X1TF U513 ( .A0(N497), .A1(N605), .B0(N488), .C0(N487), .Y(N489) );
  AOI22X1TF U514 ( .A0(XTEMP[11]), .A1(N89), .B0(SUM_AB[10]), .B1(N127), .Y(
        N488) );
  AOI21X1TF U515 ( .A0(SUM_AB[10]), .A1(N483), .B0(N496), .Y(N1001) );
  AOI22X1TF U516 ( .A0(N191), .A1(N145), .B0(N776), .B1(N775), .Y(N686) );
  AOI211X1TF U517 ( .A0(DIVISION_REMA[7]), .A1(N731), .B0(N774), .C0(N773), 
        .Y(N776) );
  OAI211X1TF U518 ( .A0(N167), .A1(N772), .B0(N771), .C0(N770), .Y(N773) );
  AOI22X1TF U519 ( .A0(N769), .A1(N768), .B0(N995), .B1(N792), .Y(N770) );
  AOI21X1TF U520 ( .A0(SUM_AB[8]), .A1(N459), .B0(N474), .Y(N995) );
  AOI32X1TF U521 ( .A0(N767), .A1(N766), .A2(N765), .B0(N764), .B1(N766), .Y(
        N768) );
  OAI32X1TF U522 ( .A0(N763), .A1(N762), .A2(X_IN[0]), .B0(N761), .B1(N763), 
        .Y(N766) );
  AOI22X1TF U523 ( .A0(DIVISION_REMA[8]), .A1(N758), .B0(SUM_AB[8]), .B1(N136), 
        .Y(N771) );
  AOI22X1TF U524 ( .A0(N472), .A1(N144), .B0(N438), .B1(N457), .Y(N714) );
  AOI21X1TF U525 ( .A0(DIVISION_HEAD[8]), .A1(N126), .B0(N431), .Y(N432) );
  OAI22X1TF U526 ( .A0(N144), .A1(N451), .B0(N504), .B1(N988), .Y(N431) );
  AOI22X1TF U527 ( .A0(DIVISION_HEAD[10]), .A1(N88), .B0(X_IN[10]), .B1(N99), 
        .Y(N434) );
  OAI22X1TF U528 ( .A0(N439), .A1(N605), .B0(N555), .B1(N473), .Y(N437) );
  OAI211X1TF U529 ( .A0(N1007), .A1(N1006), .B0(N1005), .C0(N1004), .Y(N658)
         );
  AOI22X1TF U530 ( .A0(DIVISION_HEAD[11]), .A1(N138), .B0(ZTEMP[11]), .B1(N117), .Y(N1005) );
  AOI32X1TF U531 ( .A0(N419), .A1(N457), .A2(N418), .B0(N472), .B1(N143), .Y(
        N716) );
  AOI211X1TF U532 ( .A0(DIVISION_HEAD[8]), .A1(N89), .B0(N417), .C0(N416), .Y(
        N418) );
  OAI211X1TF U533 ( .A0(N555), .A1(N449), .B0(N415), .C0(N414), .Y(N416) );
  AOI21X1TF U534 ( .A0(DIVISION_HEAD[6]), .A1(N731), .B0(N413), .Y(N414) );
  OAI22X1TF U535 ( .A0(N143), .A1(N451), .B0(N504), .B1(N982), .Y(N413) );
  OAI21X1TF U536 ( .A0(N499), .A1(N744), .B0(N410), .Y(N417) );
  AOI22X1TF U537 ( .A0(X_IN[8]), .A1(N100), .B0(X_IN[9]), .B1(N132), .Y(N410)
         );
  OAI21X1TF U538 ( .A0(N756), .A1(N178), .B0(N559), .Y(N705) );
  OAI22X1TF U539 ( .A0(N558), .A1(N557), .B0(N758), .B1(N775), .Y(N559) );
  AOI22X1TF U540 ( .A0(Y_IN[0]), .A1(N786), .B0(DIVISION_REMA[1]), .B1(N113), 
        .Y(N556) );
  AOI21X1TF U541 ( .A0(N112), .A1(N646), .B0(N973), .Y(N558) );
  INVX2TF U542 ( .A(SUM_AB[0]), .Y(N973) );
  OAI22X1TF U543 ( .A0(N191), .A1(N650), .B0(N756), .B1(N158), .Y(N693) );
  AOI21X1TF U544 ( .A0(SUM_AB[1]), .A1(N137), .B0(N649), .Y(N650) );
  AOI22X1TF U545 ( .A0(DIVISION_REMA[0]), .A1(N731), .B0(N792), .B1(N974), .Y(
        N647) );
  AOI21X1TF U546 ( .A0(SUM_AB[1]), .A1(SUM_AB[0]), .B0(N401), .Y(N974) );
  AOI22X1TF U547 ( .A0(Y_IN[1]), .A1(N786), .B0(DIVISION_REMA[2]), .B1(N114), 
        .Y(N648) );
  OAI22X1TF U548 ( .A0(N191), .A1(N748), .B0(N756), .B1(N173), .Y(N688) );
  AOI211X1TF U549 ( .A0(N989), .A1(N792), .B0(N747), .C0(N746), .Y(N748) );
  OAI211X1TF U550 ( .A0(N745), .A1(N744), .B0(N752), .C0(N743), .Y(N746) );
  AOI22X1TF U551 ( .A0(DIVISION_REMA[7]), .A1(N113), .B0(SUM_AB[6]), .B1(N136), 
        .Y(N743) );
  INVX2TF U552 ( .A(N802), .Y(N744) );
  OAI21X1TF U553 ( .A0(N200), .A1(N96), .B0(N741), .Y(N747) );
  AOI22X1TF U554 ( .A0(Y_IN[6]), .A1(N786), .B0(DIVISION_REMA[5]), .B1(N731), 
        .Y(N741) );
  AOI21X1TF U555 ( .A0(SUM_AB[6]), .A1(N440), .B0(N450), .Y(N989) );
  OAI22X1TF U556 ( .A0(N191), .A1(N736), .B0(N756), .B1(N168), .Y(N690) );
  AOI211X1TF U557 ( .A0(SUM_AB[4]), .A1(N137), .B0(N735), .C0(N734), .Y(N736)
         );
  OAI211X1TF U558 ( .A0(N733), .A1(N96), .B0(N752), .C0(N732), .Y(N734) );
  AOI22X1TF U559 ( .A0(DIVISION_REMA[5]), .A1(N114), .B0(N792), .B1(N983), .Y(
        N732) );
  AOI21X1TF U560 ( .A0(SUM_AB[4]), .A1(N420), .B0(N430), .Y(N983) );
  OAI22X1TF U561 ( .A0(N200), .A1(N799), .B0(N164), .B1(N94), .Y(N735) );
  OAI22X1TF U562 ( .A0(N191), .A1(N655), .B0(N756), .B1(N171), .Y(N692) );
  AOI211X1TF U563 ( .A0(SUM_AB[2]), .A1(N137), .B0(N654), .C0(N653), .Y(N655)
         );
  OAI211X1TF U564 ( .A0(N652), .A1(N96), .B0(N752), .C0(N651), .Y(N653) );
  AOI22X1TF U565 ( .A0(DIVISION_REMA[3]), .A1(N114), .B0(N792), .B1(N977), .Y(
        N651) );
  AOI21X1TF U566 ( .A0(SUM_AB[2]), .A1(N402), .B0(N412), .Y(N977) );
  NOR2X1TF U567 ( .A(SUM_AB[0]), .B(SUM_AB[1]), .Y(N401) );
  OAI22X1TF U568 ( .A0(N733), .A1(N799), .B0(N158), .B1(N94), .Y(N654) );
  INVX2TF U569 ( .A(N917), .Y(N906) );
  OAI211X1TF U570 ( .A0(N1016), .A1(N1015), .B0(N1014), .C0(N1013), .Y(N657)
         );
  AOI32X1TF U571 ( .A0(N1015), .A1(N1012), .A2(N1011), .B0(N1010), .B1(N1012), 
        .Y(N1013) );
  AOI211X4TF U572 ( .A0(N972), .A1(N971), .B0(N970), .C0(N116), .Y(N1012) );
  INVX2TF U573 ( .A(N966), .Y(N970) );
  AOI22X1TF U574 ( .A0(DIVISION_HEAD[12]), .A1(N138), .B0(ZTEMP[12]), .B1(N117), .Y(N1014) );
  OAI31X1TF U575 ( .A0(N964), .A1(N56), .A2(N968), .B0(N963), .Y(N965) );
  AOI31X1TF U576 ( .A0(N177), .A1(N56), .A2(N962), .B0(N961), .Y(N963) );
  AOI31X1TF U577 ( .A0(N957), .A1(N956), .A2(N955), .B0(N954), .Y(N960) );
  OAI31X1TF U578 ( .A0(N953), .A1(N952), .A2(N951), .B0(N950), .Y(N954) );
  OAI22X1TF U579 ( .A0(N510), .A1(N360), .B0(N359), .B1(N170), .Y(N723) );
  AOI211X1TF U580 ( .A0(N490), .A1(N1010), .B0(N357), .C0(N356), .Y(N360) );
  OAI31X1TF U581 ( .A0(XTEMP[12]), .A1(N358), .A2(N506), .B0(N355), .Y(N356)
         );
  INVX2TF U582 ( .A(N605), .Y(N441) );
  OAI22X1TF U583 ( .A0(N112), .A1(N1015), .B0(N499), .B1(N96), .Y(N357) );
  OAI22X1TF U584 ( .A0(N510), .A1(N509), .B0(N508), .B1(N154), .Y(N708) );
  OAI21X1TF U585 ( .A0(N504), .A1(N1006), .B0(N503), .Y(N505) );
  AOI211X1TF U586 ( .A0(SUM_AB[11]), .A1(N127), .B0(N501), .C0(N500), .Y(N503)
         );
  NAND2X2TF U587 ( .A(MODE_TYPE[1]), .B(N354), .Y(N605) );
  OAI22X1TF U588 ( .A0(N146), .A1(N93), .B0(N497), .B1(N95), .Y(N501) );
  INVX2TF U589 ( .A(N490), .Y(N504) );
  NOR2X2TF U590 ( .A(N391), .B(N1015), .Y(N490) );
  INVX2TF U591 ( .A(INTADD_0_N1), .Y(N461) );
  NOR2X1TF U592 ( .A(N151), .B(N745), .Y(INTADD_0_CI) );
  INVX2TF U593 ( .A(X_IN[0]), .Y(N745) );
  AOI31X1TF U594 ( .A0(N943), .A1(N73), .A2(N560), .B0(N351), .Y(N382) );
  OAI211X1TF U595 ( .A0(N73), .A1(N376), .B0(N361), .C0(N350), .Y(N351) );
  OAI211X1TF U596 ( .A0(N957), .A1(N349), .B0(N563), .C0(N597), .Y(N350) );
  NOR2X1TF U597 ( .A(PRE_WORK), .B(N366), .Y(N599) );
  INVX2TF U598 ( .A(N596), .Y(N563) );
  NOR2X1TF U599 ( .A(N373), .B(N945), .Y(N361) );
  INVX2TF U600 ( .A(N391), .Y(N373) );
  INVX2TF U601 ( .A(N614), .Y(N376) );
  OAI21X1TF U602 ( .A0(N756), .A1(N166), .B0(N755), .Y(N687) );
  OAI21X1TF U603 ( .A0(N754), .A1(N753), .B0(N775), .Y(N755) );
  INVX2TF U604 ( .A(N191), .Y(N775) );
  OAI211X1TF U605 ( .A0(N145), .A1(N772), .B0(N752), .C0(N751), .Y(N753) );
  AOI22X1TF U606 ( .A0(DIVISION_REMA[6]), .A1(N731), .B0(SUM_AB[7]), .B1(N136), 
        .Y(N751) );
  OAI211X1TF U607 ( .A0(N805), .A1(N994), .B0(N750), .C0(N749), .Y(N754) );
  AOI22X1TF U608 ( .A0(X_IN[1]), .A1(N802), .B0(X_IN[0]), .B1(N132), .Y(N749)
         );
  OAI21X1TF U609 ( .A0(N450), .A1(N449), .B0(N459), .Y(N994) );
  OAI22X1TF U610 ( .A0(N191), .A1(N740), .B0(N756), .B1(N165), .Y(N689) );
  AOI211X1TF U611 ( .A0(SUM_AB[5]), .A1(N137), .B0(N739), .C0(N738), .Y(N740)
         );
  OAI211X1TF U612 ( .A0(N805), .A1(N988), .B0(N752), .C0(N737), .Y(N738) );
  OAI21X1TF U613 ( .A0(N430), .A1(N429), .B0(N440), .Y(N988) );
  INVX2TF U614 ( .A(N799), .Y(N786) );
  OAI22X1TF U615 ( .A0(N191), .A1(N730), .B0(N756), .B1(N164), .Y(N691) );
  AOI211X1TF U616 ( .A0(SUM_AB[3]), .A1(N137), .B0(N729), .C0(N728), .Y(N730)
         );
  OAI211X1TF U617 ( .A0(N805), .A1(N982), .B0(N752), .C0(N727), .Y(N728) );
  AOI222X4TF U618 ( .A0(N762), .A1(N99), .B0(N760), .B1(N131), .C0(N554), .C1(
        N802), .Y(N752) );
  OAI21X1TF U619 ( .A0(N412), .A1(N411), .B0(N420), .Y(N982) );
  OAI22X1TF U620 ( .A0(N656), .A1(N799), .B0(N171), .B1(N94), .Y(N729) );
  NOR3X1TF U621 ( .A(N769), .B(N126), .C(N553), .Y(N777) );
  AOI32X1TF U622 ( .A0(N785), .A1(N811), .A2(N784), .B0(N809), .B1(N167), .Y(
        N685) );
  OAI211X1TF U623 ( .A0(N805), .A1(N1000), .B0(N781), .C0(N780), .Y(N782) );
  AOI22X1TF U624 ( .A0(DIVISION_HEAD[1]), .A1(N114), .B0(X_IN[1]), .B1(N99), 
        .Y(N780) );
  OAI21X1TF U625 ( .A0(N474), .A1(N473), .B0(N483), .Y(N1000) );
  OAI21X1TF U626 ( .A0(N779), .A1(N799), .B0(N778), .Y(N783) );
  AOI22X1TF U627 ( .A0(DIVISION_REMA[8]), .A1(N126), .B0(N795), .B1(SUM_AB[0]), 
        .Y(N778) );
  AOI22X1TF U628 ( .A0(DIVISION_HEAD[0]), .A1(N801), .B0(SUM_AB[9]), .B1(N137), 
        .Y(N785) );
  OAI21X1TF U629 ( .A0(N809), .A1(N552), .B0(N551), .Y(N706) );
  OAI21X1TF U630 ( .A0(N809), .A1(N801), .B0(DIVISION_HEAD[3]), .Y(N551) );
  AOI211X1TF U631 ( .A0(DIVISION_HEAD[2]), .A1(N126), .B0(N550), .C0(N549), 
        .Y(N552) );
  AOI22X1TF U632 ( .A0(N795), .A1(SUM_AB[3]), .B0(N1010), .B1(N792), .Y(N546)
         );
  NOR2X1TF U633 ( .A(N1015), .B(N1011), .Y(N1010) );
  AOI22X1TF U634 ( .A0(N943), .A1(SUM_AB[12]), .B0(X_IN[5]), .B1(N132), .Y(
        N547) );
  AOI22X1TF U635 ( .A0(X_IN[4]), .A1(N100), .B0(X_IN[6]), .B1(N802), .Y(N548)
         );
  OAI22X1TF U636 ( .A0(N545), .A1(N799), .B0(N544), .B1(N96), .Y(N550) );
  AOI32X1TF U637 ( .A0(N812), .A1(N811), .A2(N810), .B0(N809), .B1(N161), .Y(
        N683) );
  AOI211X1TF U638 ( .A0(DIVISION_HEAD[3]), .A1(N114), .B0(N807), .C0(N806), 
        .Y(N810) );
  OAI211X1TF U639 ( .A0(N805), .A1(N1006), .B0(N804), .C0(N803), .Y(N806) );
  AOI22X1TF U640 ( .A0(X_IN[3]), .A1(N99), .B0(X_IN[5]), .B1(N802), .Y(N803)
         );
  AND2X2TF U641 ( .A(N759), .B(N764), .Y(N761) );
  INVX2TF U642 ( .A(N383), .Y(N769) );
  AOI22X1TF U643 ( .A0(DIVISION_HEAD[1]), .A1(N126), .B0(DIVISION_HEAD[2]), 
        .B1(N801), .Y(N804) );
  INVX2TF U644 ( .A(N451), .Y(N801) );
  OAI21X1TF U645 ( .A0(N496), .A1(N495), .B0(N1011), .Y(N1006) );
  INVX2TF U646 ( .A(SUM_AB[11]), .Y(N495) );
  INVX2TF U647 ( .A(SUM_AB[9]), .Y(N473) );
  INVX2TF U648 ( .A(SUM_AB[7]), .Y(N449) );
  NOR2X1TF U649 ( .A(SUM_AB[6]), .B(N440), .Y(N450) );
  INVX2TF U650 ( .A(SUM_AB[5]), .Y(N429) );
  NOR2X1TF U651 ( .A(SUM_AB[4]), .B(N420), .Y(N430) );
  INVX2TF U652 ( .A(SUM_AB[3]), .Y(N411) );
  NOR3X1TF U653 ( .A(SUM_AB[0]), .B(SUM_AB[2]), .C(SUM_AB[1]), .Y(N412) );
  INVX2TF U654 ( .A(N792), .Y(N805) );
  NOR2X2TF U655 ( .A(N1015), .B(N646), .Y(N792) );
  INVX2TF U656 ( .A(SUM_AB[12]), .Y(N1015) );
  OAI21X1TF U657 ( .A0(N800), .A1(N799), .B0(N798), .Y(N807) );
  INVX2TF U658 ( .A(N95), .Y(N797) );
  NAND2X2TF U659 ( .A(N354), .B(N313), .Y(N799) );
  INVX2TF U660 ( .A(N809), .Y(N811) );
  INVX2TF U661 ( .A(N354), .Y(N636) );
  AOI31X1TF U662 ( .A0(N122), .A1(N381), .A2(N380), .B0(N379), .Y(N543) );
  INVX2TF U663 ( .A(N306), .Y(N760) );
  OAI211X1TF U664 ( .A0(X_IN[12]), .A1(N544), .B0(N305), .C0(N304), .Y(N306)
         );
  OAI22X1TF U665 ( .A0(Y_IN[10]), .A1(N303), .B0(N302), .B1(N301), .Y(N304) );
  OAI22X1TF U666 ( .A0(X_IN[10]), .A1(N300), .B0(X_IN[11]), .B1(N779), .Y(N301) );
  OAI21X1TF U667 ( .A0(Y_IN[9]), .A1(N299), .B0(Y_IN[8]), .Y(N300) );
  AOI211X1TF U668 ( .A0(X_IN[10]), .A1(N757), .B0(N298), .C0(N297), .Y(N302)
         );
  AOI21X1TF U669 ( .A0(Y_IN[7]), .A1(N497), .B0(N296), .Y(N297) );
  AOI211X1TF U670 ( .A0(X_IN[8]), .A1(N295), .B0(N294), .C0(N293), .Y(N296) );
  NOR2X1TF U671 ( .A(N84), .B(N497), .Y(N294) );
  AOI21X1TF U672 ( .A0(N192), .A1(N465), .B0(N292), .Y(N295) );
  AOI211X1TF U673 ( .A0(X_IN[6]), .A1(N291), .B0(N290), .C0(N289), .Y(N292) );
  NOR2X1TF U674 ( .A(N192), .B(N465), .Y(N290) );
  AOI32X1TF U675 ( .A0(N288), .A1(N287), .A2(N317), .B0(N286), .B1(N287), .Y(
        N291) );
  OAI22X1TF U676 ( .A0(X_IN[4]), .A1(N733), .B0(N101), .B1(N656), .Y(N286) );
  OAI32X1TF U677 ( .A0(N285), .A1(N85), .A2(N315), .B0(X_IN[2]), .B1(N285), 
        .Y(N288) );
  INVX2TF U678 ( .A(X_IN[7]), .Y(N465) );
  INVX2TF U679 ( .A(X_IN[9]), .Y(N497) );
  NOR2X1TF U680 ( .A(Y_IN[9]), .B(N299), .Y(N298) );
  INVX2TF U681 ( .A(X_IN[11]), .Y(N299) );
  NOR2X1TF U682 ( .A(Y_IN[12]), .B(Y_IN[11]), .Y(N305) );
  INVX2TF U683 ( .A(N765), .Y(N554) );
  OR2X2TF U684 ( .A(MODE_TYPE[0]), .B(N313), .Y(N764) );
  INVX2TF U685 ( .A(MODE_TYPE[1]), .Y(N313) );
  OAI31X1TF U686 ( .A0(N281), .A1(N280), .A2(N279), .B0(N278), .Y(N282) );
  NOR2X1TF U687 ( .A(X_IN[10]), .B(N779), .Y(N279) );
  AOI211X1TF U688 ( .A0(X_IN[10]), .A1(N779), .B0(X_IN[9]), .C0(N757), .Y(N280) );
  AOI211X1TF U689 ( .A0(X_IN[9]), .A1(N757), .B0(N277), .C0(N276), .Y(N281) );
  AOI21X1TF U690 ( .A0(Y_IN[7]), .A1(N485), .B0(N275), .Y(N276) );
  AOI211X1TF U691 ( .A0(N274), .A1(X_IN[7]), .B0(N273), .C0(N272), .Y(N275) );
  NOR2X1TF U692 ( .A(Y_IN[7]), .B(N485), .Y(N273) );
  AOI21X1TF U693 ( .A0(N192), .A1(N460), .B0(N271), .Y(N274) );
  AOI211X1TF U694 ( .A0(N270), .A1(X_IN[5]), .B0(N269), .C0(N268), .Y(N271) );
  NOR2X1TF U695 ( .A(N192), .B(N460), .Y(N269) );
  AOI211X1TF U696 ( .A0(Y_IN[3]), .A1(N439), .B0(N267), .C0(N266), .Y(N270) );
  AOI211X1TF U697 ( .A0(X_IN[4]), .A1(N656), .B0(N85), .C0(N733), .Y(N266) );
  OAI32X1TF U698 ( .A0(N265), .A1(X_IN[2]), .A2(N315), .B0(X_IN[1]), .B1(N265), 
        .Y(N267) );
  OAI211X1TF U699 ( .A0(Y_IN[3]), .A1(N439), .B0(N264), .C0(N317), .Y(N265) );
  AOI22X1TF U700 ( .A0(N85), .A1(N733), .B0(X_IN[2]), .B1(N316), .Y(N264) );
  INVX2TF U701 ( .A(X_IN[4]), .Y(N439) );
  INVX2TF U702 ( .A(X_IN[6]), .Y(N460) );
  INVX2TF U703 ( .A(X_IN[8]), .Y(N485) );
  NOR2X1TF U704 ( .A(Y_IN[9]), .B(N499), .Y(N277) );
  INVX2TF U705 ( .A(X_IN[10]), .Y(N499) );
  NOR2X1TF U706 ( .A(Y_IN[11]), .B(N303), .Y(N283) );
  INVX2TF U707 ( .A(X_IN[12]), .Y(N303) );
  INVX2TF U708 ( .A(N340), .Y(N381) );
  AOI22X1TF U709 ( .A0(N795), .A1(SUM_AB[2]), .B0(SUM_AB[11]), .B1(N137), .Y(
        N812) );
  OAI21X1TF U710 ( .A0(N170), .A1(N109), .B0(N257), .Y(OPER_A[12]) );
  INVX2TF U711 ( .A(N555), .Y(N795) );
  OAI211X1TF U712 ( .A0(N857), .A1(N856), .B0(N855), .C0(N854), .Y(N678) );
  AOI32X1TF U713 ( .A0(N933), .A1(OPER_B[4]), .A2(N853), .B0(N878), .B1(
        OPER_B[4]), .Y(N854) );
  AOI211X1TF U714 ( .A0(N858), .A1(OPER_B[5]), .B0(N852), .C0(N851), .Y(N855)
         );
  OAI31X1TF U715 ( .A0(N930), .A1(OPER_A[4]), .A2(N850), .B0(N204), .Y(N851)
         );
  AOI21X1TF U716 ( .A0(N104), .A1(C152_DATA4_4), .B0(N205), .Y(N204) );
  NOR3X1TF U717 ( .A(OPER_B[4]), .B(N853), .C(N107), .Y(N852) );
  AOI21X1TF U718 ( .A0(N927), .A1(N850), .B0(N849), .Y(N856) );
  OR2X2TF U719 ( .A(N825), .B(N827), .Y(N210) );
  AOI21X1TF U720 ( .A0(N927), .A1(N826), .B0(N849), .Y(N825) );
  INVX2TF U721 ( .A(N928), .Y(N849) );
  AOI21X1TF U722 ( .A0(N105), .A1(C152_DATA4_1), .B0(N879), .Y(N211) );
  AOI211X1TF U723 ( .A0(N858), .A1(OPER_B[2]), .B0(N823), .C0(N822), .Y(N824)
         );
  NOR3X1TF U724 ( .A(N826), .B(OPER_A[1]), .C(N930), .Y(N822) );
  INVX2TF U725 ( .A(OPER_A[0]), .Y(N826) );
  OAI32X1TF U726 ( .A0(N181), .A1(OPER_B[0]), .A2(N107), .B0(N931), .B1(N181), 
        .Y(N823) );
  OAI31X1TF U727 ( .A0(OPER_B[1]), .A1(N107), .A2(N183), .B0(N820), .Y(N821)
         );
  OAI21X1TF U728 ( .A0(N152), .A1(N98), .B0(N232), .Y(FOUT[4]) );
  AOI21X1TF U729 ( .A0(N221), .A1(DIVISION_REMA[4]), .B0(N231), .Y(N232) );
  OAI22X1TF U730 ( .A0(N153), .A1(N87), .B0(N173), .B1(N81), .Y(N231) );
  OAI211X1TF U731 ( .A0(SIGN_Y), .A1(N962), .B0(N222), .C0(N968), .Y(N893) );
  INVX2TF U732 ( .A(N882), .Y(N858) );
  OAI21X1TF U733 ( .A0(N142), .A1(N97), .B0(N226), .Y(FOUT[1]) );
  AOI21X1TF U734 ( .A0(N221), .A1(DIVISION_REMA[1]), .B0(N225), .Y(N226) );
  OAI22X1TF U735 ( .A0(N143), .A1(N86), .B0(N164), .B1(N80), .Y(N225) );
  AOI22X1TF U736 ( .A0(OPER_B[9]), .A1(N901), .B0(OPER_A[9]), .B1(N900), .Y(
        N902) );
  OAI21X1TF U737 ( .A0(N930), .A1(N899), .B0(N928), .Y(N900) );
  OAI21X1TF U738 ( .A0(N107), .A1(N898), .B0(N931), .Y(N901) );
  AOI31X1TF U739 ( .A0(N933), .A1(N187), .A2(N898), .B0(N897), .Y(N903) );
  OAI211X1TF U740 ( .A0(N160), .A1(N940), .B0(N207), .C0(N206), .Y(N897) );
  AOI22X1TF U741 ( .A0(SIGN_Y), .A1(N895), .B0(N894), .B1(N899), .Y(N904) );
  NOR2X1TF U742 ( .A(N930), .B(OPER_A[9]), .Y(N894) );
  OR2X2TF U743 ( .A(N925), .B(N879), .Y(N205) );
  NOR2X1TF U744 ( .A(N964), .B(N831), .Y(N864) );
  INVX2TF U745 ( .A(N931), .Y(N878) );
  OAI211X1TF U746 ( .A0(N186), .A1(N940), .B0(N939), .C0(N938), .Y(N671) );
  AOI211X1TF U747 ( .A0(OPER_A[11]), .A1(N937), .B0(N936), .C0(N935), .Y(N938)
         );
  AOI21X1TF U748 ( .A0(N961), .A1(N222), .B0(N208), .Y(N209) );
  NOR3X1TF U749 ( .A(N106), .B(OPER_B[11]), .C(N934), .Y(N208) );
  INVX2TF U750 ( .A(N932), .Y(N934) );
  NOR3X1TF U751 ( .A(N73), .B(N177), .C(N962), .Y(N961) );
  OAI22X1TF U752 ( .A0(N189), .A1(N200), .B0(N201), .B1(OFFSET[2]), .Y(C2_Z_4)
         );
  INVX2TF U753 ( .A(Y_IN[4]), .Y(N200) );
  OAI22X1TF U754 ( .A0(N189), .A1(N199), .B0(N201), .B1(OFFSET[3]), .Y(C2_Z_5)
         );
  OAI22X1TF U755 ( .A0(N189), .A1(N198), .B0(N201), .B1(OFFSET[4]), .Y(C2_Z_6)
         );
  OAI22X1TF U756 ( .A0(N189), .A1(N193), .B0(N201), .B1(OFFSET[5]), .Y(C2_Z_7)
         );
  OAI22X1TF U757 ( .A0(N189), .A1(N757), .B0(N201), .B1(OFFSET[6]), .Y(C2_Z_8)
         );
  OAI22X1TF U758 ( .A0(N189), .A1(N779), .B0(N201), .B1(OFFSET[7]), .Y(C2_Z_9)
         );
  OAI22X1TF U759 ( .A0(N189), .A1(N544), .B0(N133), .B1(OFFSET[8]), .Y(C2_Z_10) );
  OAI22X1TF U760 ( .A0(N189), .A1(N800), .B0(N133), .B1(OFFSET[9]), .Y(C2_Z_11) );
  INVX2TF U761 ( .A(Y_IN[11]), .Y(N800) );
  OAI32X1TF U762 ( .A0(N184), .A1(N932), .A2(N107), .B0(N931), .B1(N184), .Y(
        N936) );
  NOR2X1TF U763 ( .A(OPER_B[9]), .B(N898), .Y(N918) );
  NOR2X1TF U764 ( .A(N863), .B(OPER_B[6]), .Y(N880) );
  INVX2TF U765 ( .A(N867), .Y(N863) );
  NOR2X1TF U766 ( .A(OPER_B[5]), .B(N859), .Y(N867) );
  NOR2X1TF U767 ( .A(OPER_B[3]), .B(N842), .Y(N853) );
  OAI21X1TF U768 ( .A0(N930), .A1(N929), .B0(N928), .Y(N937) );
  AOI31X1TF U769 ( .A0(N927), .A1(N926), .A2(N929), .B0(N925), .Y(N939) );
  AOI211X1TF U770 ( .A0(N56), .A1(N962), .B0(SIGN_Y), .C0(N905), .Y(N925) );
  NOR2X1TF U771 ( .A(OPER_A[9]), .B(N899), .Y(N912) );
  NOR2X1TF U772 ( .A(OPER_A[7]), .B(N881), .Y(N886) );
  NOR2X1TF U773 ( .A(OPER_A[5]), .B(N860), .Y(N870) );
  NOR2X1TF U774 ( .A(OPER_A[3]), .B(N841), .Y(N850) );
  OAI21X1TF U775 ( .A0(N152), .A1(N109), .B0(N248), .Y(OPER_A[4]) );
  OAI21X1TF U776 ( .A0(N144), .A1(N109), .B0(N249), .Y(OPER_A[5]) );
  OAI21X1TF U777 ( .A0(N153), .A1(N109), .B0(N250), .Y(OPER_A[6]) );
  OAI21X1TF U778 ( .A0(N141), .A1(N109), .B0(N251), .Y(OPER_A[7]) );
  OAI21X1TF U779 ( .A0(N175), .A1(N109), .B0(N252), .Y(OPER_A[8]) );
  OAI21X1TF U780 ( .A0(N109), .A1(N525), .B0(N253), .Y(OPER_A[9]) );
  OAI21X1TF U781 ( .A0(N109), .A1(N146), .B0(N254), .Y(OPER_A[10]) );
  OAI21X1TF U782 ( .A0(N109), .A1(N154), .B0(N255), .Y(OPER_A[11]) );
  OAI211X1TF U783 ( .A0(N176), .A1(N940), .B0(N848), .C0(N847), .Y(N679) );
  AOI211X1TF U784 ( .A0(OPER_A[3]), .A1(N846), .B0(N845), .C0(N844), .Y(N847)
         );
  OAI31X1TF U785 ( .A0(N930), .A1(OPER_A[3]), .A2(N843), .B0(N203), .Y(N844)
         );
  AOI21X1TF U786 ( .A0(C152_DATA4_3), .A1(N104), .B0(N895), .Y(N203) );
  OAI22X1TF U787 ( .A0(N967), .A1(N656), .B0(N201), .B1(OFFSET[1]), .Y(C2_Z_3)
         );
  INVX2TF U788 ( .A(DP_OP_333_124_4748_N57), .Y(N201) );
  INVX2TF U789 ( .A(Y_IN[3]), .Y(N656) );
  OAI32X1TF U790 ( .A0(N182), .A1(N106), .A2(N842), .B0(N931), .B1(N182), .Y(
        N845) );
  INVX2TF U791 ( .A(N862), .Y(N916) );
  AOI32X1TF U792 ( .A0(N602), .A1(N348), .A2(N819), .B0(N947), .B1(N347), .Y(
        N862) );
  INVX2TF U793 ( .A(N942), .Y(N947) );
  OAI21X1TF U794 ( .A0(N930), .A1(N841), .B0(N928), .Y(N846) );
  INVX2TF U795 ( .A(N832), .Y(N907) );
  AOI21X1TF U796 ( .A0(N561), .A1(N347), .B0(N560), .Y(N832) );
  INVX2TF U797 ( .A(N843), .Y(N841) );
  NOR3X1TF U798 ( .A(OPER_A[2]), .B(OPER_A[1]), .C(OPER_A[0]), .Y(N843) );
  OAI21X1TF U799 ( .A0(N150), .A1(N108), .B0(N246), .Y(OPER_A[2]) );
  INVX2TF U800 ( .A(N927), .Y(N930) );
  NOR2X2TF U801 ( .A(N919), .B(N911), .Y(N927) );
  INVX2TF U802 ( .A(N892), .Y(N919) );
  OAI21X1TF U803 ( .A0(N143), .A1(N108), .B0(N247), .Y(OPER_A[3]) );
  AOI31X1TF U804 ( .A0(N933), .A1(N182), .A2(N842), .B0(N876), .Y(N848) );
  OAI21X1TF U805 ( .A0(N972), .A1(N905), .B0(N838), .Y(N876) );
  INVX2TF U806 ( .A(N905), .Y(N222) );
  INVX2TF U807 ( .A(N346), .Y(N956) );
  INVX2TF U808 ( .A(N562), .Y(N949) );
  NOR2X1TF U809 ( .A(OPER_B[1]), .B(OPER_B[0]), .Y(N834) );
  INVX2TF U810 ( .A(N347), .Y(N348) );
  INVX2TF U811 ( .A(N602), .Y(N818) );
  NOR2X2TF U812 ( .A(N600), .B(N628), .Y(N819) );
  AOI221X1TF U813 ( .A0(N128), .A1(N157), .B0(N180), .B1(N91), .C0(N814), .Y(
        N815) );
  AOI22X1TF U814 ( .A0(\INDEX[2] ), .A1(N90), .B0(N124), .B1(\RSHT_BITS[3] ), 
        .Y(N813) );
  AOI32X1TF U815 ( .A0(N942), .A1(N950), .A2(N370), .B0(N952), .B1(N950), .Y(
        N344) );
  OR2X2TF U816 ( .A(N628), .B(N148), .Y(N370) );
  INVX2TF U817 ( .A(N600), .Y(N639) );
  OAI21X1TF U818 ( .A0(N346), .A1(N941), .B0(N342), .Y(N604) );
  OAI21X1TF U819 ( .A0(N567), .A1(N561), .B0(N343), .Y(N342) );
  NOR2X2TF U820 ( .A(\RSHT_BITS[3] ), .B(N588), .Y(N602) );
  NOR3X1TF U821 ( .A(N121), .B(N122), .C(N951), .Y(N817) );
  INVX2TF U822 ( .A(N957), .Y(N964) );
  NOR2X1TF U823 ( .A(SIGN_Y), .B(N110), .Y(N896) );
  INVX2TF U824 ( .A(N310), .Y(N624) );
  OAI22X1TF U825 ( .A0(Y_IN[12]), .A1(N175), .B0(N338), .B1(N337), .Y(N339) );
  OAI31X1TF U826 ( .A0(N336), .A1(DIVISION_HEAD[10]), .A2(N544), .B0(N335), 
        .Y(N337) );
  AOI22X1TF U827 ( .A0(Y_IN[11]), .A1(N141), .B0(N334), .B1(N333), .Y(N335) );
  OAI22X1TF U828 ( .A0(DIVISION_HEAD[8]), .A1(N757), .B0(DIVISION_HEAD[9]), 
        .B1(N779), .Y(N333) );
  INVX2TF U829 ( .A(N332), .Y(N334) );
  NOR2X1TF U830 ( .A(Y_IN[11]), .B(N141), .Y(N336) );
  AOI211X1TF U831 ( .A0(DIVISION_HEAD[8]), .A1(N757), .B0(N331), .C0(N332), 
        .Y(N338) );
  OAI21X1TF U832 ( .A0(Y_IN[11]), .A1(N141), .B0(N330), .Y(N332) );
  AOI22X1TF U833 ( .A0(DIVISION_HEAD[10]), .A1(N544), .B0(DIVISION_HEAD[9]), 
        .B1(N779), .Y(N330) );
  INVX2TF U834 ( .A(Y_IN[9]), .Y(N779) );
  INVX2TF U835 ( .A(Y_IN[10]), .Y(N544) );
  AOI21X1TF U836 ( .A0(N84), .A1(N143), .B0(N329), .Y(N331) );
  AOI211X1TF U837 ( .A0(N328), .A1(DIVISION_HEAD[6]), .B0(N327), .C0(N326), 
        .Y(N329) );
  NOR2X1TF U838 ( .A(N84), .B(N143), .Y(N327) );
  AOI21X1TF U839 ( .A0(N192), .A1(N142), .B0(N325), .Y(N328) );
  AOI211X1TF U840 ( .A0(N324), .A1(DIVISION_HEAD[4]), .B0(N323), .C0(N322), 
        .Y(N325) );
  NOR2X1TF U841 ( .A(Y_IN[5]), .B(N142), .Y(N323) );
  AOI21X1TF U842 ( .A0(Y_IN[3]), .A1(N147), .B0(N321), .Y(N324) );
  OAI32X1TF U843 ( .A0(N320), .A1(DIVISION_HEAD[2]), .A2(N733), .B0(N319), 
        .B1(N320), .Y(N321) );
  OAI211X1TF U844 ( .A0(Y_IN[2]), .A1(N161), .B0(N318), .C0(N317), .Y(N319) );
  INVX2TF U845 ( .A(Y_IN[0]), .Y(N652) );
  INVX2TF U846 ( .A(Y_IN[1]), .Y(N315) );
  INVX2TF U847 ( .A(Y_IN[2]), .Y(N733) );
  NOR2X1TF U848 ( .A(Y_IN[3]), .B(N147), .Y(N320) );
  INVX2TF U849 ( .A(Y_IN[8]), .Y(N757) );
  INVX2TF U850 ( .A(Y_IN[12]), .Y(N545) );
  OAI21X1TF U851 ( .A0(N175), .A1(N98), .B0(N240), .Y(FOUT[8]) );
  AOI21X1TF U852 ( .A0(N221), .A1(DIVISION_REMA[8]), .B0(N239), .Y(N240) );
  OAI22X1TF U853 ( .A0(N172), .A1(N81), .B0(N146), .B1(N86), .Y(N239) );
  OAI21X1TF U854 ( .A0(N144), .A1(N97), .B0(N234), .Y(FOUT[5]) );
  AOI21X1TF U855 ( .A0(N221), .A1(DIVISION_REMA[5]), .B0(N233), .Y(N234) );
  OAI22X1TF U856 ( .A0(N141), .A1(N86), .B0(N166), .B1(N80), .Y(N233) );
  OAI21X1TF U857 ( .A0(N141), .A1(N98), .B0(N238), .Y(FOUT[7]) );
  AOI21X1TF U858 ( .A0(N221), .A1(DIVISION_REMA[7]), .B0(N237), .Y(N238) );
  OAI22X1TF U859 ( .A0(N167), .A1(N81), .B0(N525), .B1(N87), .Y(N237) );
  OAI21X1TF U860 ( .A0(N143), .A1(N97), .B0(N230), .Y(FOUT[3]) );
  AOI21X1TF U861 ( .A0(N221), .A1(DIVISION_REMA[3]), .B0(N229), .Y(N230) );
  OAI22X1TF U862 ( .A0(N144), .A1(N86), .B0(N165), .B1(N80), .Y(N229) );
  OAI21X1TF U863 ( .A0(N153), .A1(N98), .B0(N236), .Y(FOUT[6]) );
  AOI21X1TF U864 ( .A0(N221), .A1(DIVISION_REMA[6]), .B0(N235), .Y(N236) );
  OAI22X1TF U865 ( .A0(N175), .A1(N87), .B0(N145), .B1(N80), .Y(N235) );
  OAI21X1TF U866 ( .A0(N150), .A1(N97), .B0(N228), .Y(FOUT[2]) );
  AOI21X1TF U867 ( .A0(N221), .A1(DIVISION_REMA[2]), .B0(N227), .Y(N228) );
  OAI22X1TF U868 ( .A0(N152), .A1(N86), .B0(N168), .B1(N80), .Y(N227) );
  NOR2X1TF U869 ( .A(N340), .B(N371), .Y(ALU_IS_DONE) );
  OAI211X1TF U870 ( .A0(N150), .A1(N87), .B0(N224), .C0(N223), .Y(FOUT[0]) );
  AOI22X1TF U871 ( .A0(N119), .A1(\INTADD_0_SUM[5] ), .B0(N795), .B1(
        SUM_AB[10]), .Y(N445) );
  AOI21X1TF U872 ( .A0(N119), .A1(N469), .B0(N468), .Y(N470) );
  AOI22X1TF U873 ( .A0(N118), .A1(N462), .B0(SUM_AB[8]), .B1(N127), .Y(N464)
         );
  AOI31X1TF U874 ( .A0(X_IN[0]), .A1(N119), .A2(N151), .B0(N387), .Y(N388) );
  AOI22X1TF U875 ( .A0(N119), .A1(\INTADD_0_SUM[1] ), .B0(SUM_AB[2]), .B1(N130), .Y(N409) );
  AOI22X1TF U876 ( .A0(N119), .A1(\INTADD_0_SUM[3] ), .B0(SUM_AB[4]), .B1(N130), .Y(N428) );
  AOI22X1TF U877 ( .A0(N119), .A1(\INTADD_0_SUM[0] ), .B0(SUM_AB[1]), .B1(N130), .Y(N399) );
  AOI22X1TF U878 ( .A0(N119), .A1(\INTADD_0_SUM[6] ), .B0(SUM_AB[7]), .B1(N130), .Y(N458) );
  AOI31X1TF U879 ( .A0(N118), .A1(N146), .A2(N491), .B0(N486), .Y(N487) );
  AOI22X1TF U880 ( .A0(N118), .A1(\INTADD_0_SUM[4] ), .B0(SUM_AB[5]), .B1(N127), .Y(N435) );
  AOI22X1TF U881 ( .A0(N119), .A1(\INTADD_0_SUM[2] ), .B0(SUM_AB[3]), .B1(N130), .Y(N419) );
  AOI21X1TF U882 ( .A0(N119), .A1(N358), .B0(N510), .Y(N359) );
  AOI31X1TF U883 ( .A0(N119), .A1(N154), .A2(N507), .B0(N505), .Y(N509) );
  NOR2X1TF U884 ( .A(ALU_TYPE[2]), .B(ALU_TYPE[0]), .Y(N196) );
  NAND3X1TF U885 ( .A(N893), .B(N216), .C(N215), .Y(N674) );
  NAND4BX1TF U886 ( .AN(N839), .B(N213), .C(N840), .D(N212), .Y(N680) );
  AOI2BB2X1TF U887 ( .B0(N105), .B1(C152_DATA4_2), .A0N(N155), .A1N(N924), .Y(
        N212) );
  OAI2BB1X1TF U888 ( .A0N(N105), .A1N(C152_DATA4_10), .B0(N217), .Y(N672) );
  NAND4BX1TF U889 ( .AN(N821), .B(N824), .C(N211), .D(N210), .Y(N681) );
  OR3X1TF U890 ( .A(N905), .B(N74), .C(N896), .Y(N206) );
  NAND2X1TF U891 ( .A(N104), .B(C152_DATA4_9), .Y(N207) );
  OAI2BB1X1TF U892 ( .A0N(N104), .A1N(C152_DATA4_11), .B0(N209), .Y(N935) );
  OAI2BB2XLTF U893 ( .B0(OFFSET[0]), .B1(N201), .A0N(Y_IN[2]), .A1N(N125), .Y(
        C2_Z_2) );
  AOI2BB2X1TF U894 ( .B0(N221), .B1(DIVISION_REMA[0]), .A0N(N171), .A1N(N81), 
        .Y(N224) );
  OAI222X1TF U895 ( .A0(N97), .A1(N525), .B0(N81), .B1(N161), .C0(N154), .C1(
        N87), .Y(FOUT[9]) );
  NAND2X1TF U896 ( .A(N148), .B(N163), .Y(N371) );
  NAND3X1TF U897 ( .A(STEP[2]), .B(STEP[3]), .C(N639), .Y(N942) );
  NAND3X1TF U898 ( .A(N542), .B(N383), .C(N631), .Y(N644) );
  NOR4XLTF U899 ( .A(N758), .B(N614), .C(N797), .D(N644), .Y(N263) );
  AOI222XLTF U900 ( .A0(STEP[2]), .A1(N149), .B0(N121), .B1(N163), .C0(N140), 
        .C1(N122), .Y(N261) );
  NAND3X1TF U901 ( .A(N263), .B(N362), .C(N630), .Y(N616) );
  AOI2BB1X1TF U902 ( .A0N(X_IN[5]), .A1N(N270), .B0(Y_IN[4]), .Y(N268) );
  AOI2BB1X1TF U903 ( .A0N(X_IN[7]), .A1N(N274), .B0(Y_IN[6]), .Y(N272) );
  NAND2X1TF U904 ( .A(MODE_TYPE[0]), .B(N313), .Y(N759) );
  AO22X1TF U905 ( .A0(X_IN[4]), .A1(N733), .B0(N85), .B1(N316), .Y(N285) );
  NAND2X1TF U906 ( .A(N101), .B(N656), .Y(N287) );
  AOI2BB1X1TF U907 ( .A0N(N291), .A1N(X_IN[6]), .B0(Y_IN[4]), .Y(N289) );
  AOI2BB1X1TF U908 ( .A0N(N295), .A1N(X_IN[8]), .B0(Y_IN[6]), .Y(N293) );
  NAND2X1TF U909 ( .A(N156), .B(N180), .Y(N613) );
  NAND4BX1TF U910 ( .AN(N379), .B(N314), .C(N799), .D(N362), .Y(N725) );
  NAND2X1TF U911 ( .A(N834), .B(N155), .Y(N842) );
  NAND2X1TF U912 ( .A(N853), .B(N176), .Y(N859) );
  NOR2BX1TF U913 ( .AN(N880), .B(OPER_B[7]), .Y(N883) );
  NAND2X1TF U914 ( .A(N883), .B(N159), .Y(N898) );
  NAND2X1TF U915 ( .A(N918), .B(N160), .Y(N932) );
  NAND2X1TF U916 ( .A(N896), .B(N74), .Y(N955) );
  NAND2X1TF U917 ( .A(N562), .B(N955), .Y(N941) );
  NAND2X1TF U918 ( .A(N964), .B(N377), .Y(N570) );
  NAND3X1TF U919 ( .A(N92), .B(N91), .C(N90), .Y(N588) );
  NOR2BX1TF U920 ( .AN(N570), .B(N602), .Y(N567) );
  NAND2X1TF U921 ( .A(PRE_WORK), .B(N352), .Y(N950) );
  NAND2X1TF U922 ( .A(N602), .B(N819), .Y(N345) );
  NAND2X1TF U923 ( .A(N220), .B(N956), .Y(N364) );
  NAND3X1TF U924 ( .A(SIGN_Y), .B(N74), .C(N895), .Y(N820) );
  NAND2X1TF U925 ( .A(N857), .B(N850), .Y(N860) );
  NAND2X1TF U926 ( .A(N869), .B(N870), .Y(N881) );
  NAND2X1TF U927 ( .A(N885), .B(N886), .Y(N899) );
  NAND2X1TF U928 ( .A(N910), .B(N912), .Y(N929) );
  NAND3X1TF U929 ( .A(N602), .B(N599), .C(N162), .Y(N597) );
  NAND2X1TF U930 ( .A(N412), .B(N411), .Y(N420) );
  NAND2X1TF U931 ( .A(N430), .B(N429), .Y(N440) );
  NAND2X1TF U932 ( .A(N450), .B(N449), .Y(N459) );
  NAND2X1TF U933 ( .A(N496), .B(N495), .Y(N1011) );
  AOI222XLTF U934 ( .A0(XTEMP[11]), .A1(X_IN[11]), .B0(XTEMP[11]), .B1(N494), 
        .C0(X_IN[11]), .C1(N494), .Y(N353) );
  XOR2X1TF U935 ( .A(X_IN[12]), .B(N353), .Y(N358) );
  NAND3X1TF U936 ( .A(N563), .B(POST_WORK), .C(N599), .Y(N374) );
  NAND3BX1TF U937 ( .AN(N364), .B(N949), .C(N964), .Y(N595) );
  NAND3X1TF U938 ( .A(N606), .B(N365), .C(N595), .Y(N944) );
  NAND2X1TF U939 ( .A(N112), .B(N391), .Y(N378) );
  NAND3X1TF U940 ( .A(N381), .B(N122), .C(DP_OP_333_124_4748_N57), .Y(N635) );
  NOR2BX1TF U941 ( .AN(N631), .B(N945), .Y(N539) );
  NAND4X1TF U942 ( .A(N424), .B(N423), .C(N422), .D(N421), .Y(N425) );
  NAND4X1TF U943 ( .A(N435), .B(N434), .C(N433), .D(N432), .Y(N436) );
  NAND4X1TF U944 ( .A(N445), .B(N444), .C(N443), .D(N442), .Y(N446) );
  OAI2BB1X1TF U945 ( .A0N(DIVISION_HEAD[10]), .A1N(N468), .B0(N448), .Y(N713)
         );
  AOI2BB2X1TF U946 ( .B0(X_IN[9]), .B1(N475), .A0N(N475), .A1N(X_IN[9]), .Y(
        N480) );
  NAND3X1TF U947 ( .A(N118), .B(N525), .C(N480), .Y(N476) );
  AOI2BB1X1TF U948 ( .A0N(N506), .A1N(N480), .B0(N510), .Y(N481) );
  AOI2BB2X1TF U949 ( .B0(N484), .B1(N499), .A0N(N499), .A1N(N484), .Y(N491) );
  AOI2BB1X1TF U950 ( .A0N(N506), .A1N(N491), .B0(N510), .Y(N492) );
  AOI2BB2X1TF U951 ( .B0(N79), .B1(N494), .A0N(N494), .A1N(N79), .Y(N507) );
  OAI2BB2XLTF U952 ( .B0(N499), .B1(N605), .A0N(XTEMP[12]), .A1N(N88), .Y(N500) );
  AOI2BB1X1TF U953 ( .A0N(N506), .A1N(N507), .B0(N510), .Y(N508) );
  AOI2BB1X1TF U954 ( .A0N(DIVISION_REMA[2]), .A1N(N514), .B0(DIVISION_HEAD[6]), 
        .Y(N512) );
  OA21XLTF U955 ( .A0(N152), .A1(DIVISION_REMA[4]), .B0(N516), .Y(N518) );
  OA21XLTF U956 ( .A0(N153), .A1(DIVISION_REMA[6]), .B0(N520), .Y(N522) );
  OA21XLTF U957 ( .A0(XTEMP[12]), .A1(N532), .B0(N147), .Y(N531) );
  NAND4X1TF U958 ( .A(N542), .B(N541), .C(N635), .D(N540), .Y(N553) );
  NAND3X1TF U959 ( .A(N548), .B(N547), .C(N546), .Y(N549) );
  NAND3X1TF U960 ( .A(N752), .B(N556), .C(N555), .Y(N557) );
  NAND3X1TF U961 ( .A(N563), .B(N599), .C(N818), .Y(N569) );
  NAND4X1TF U962 ( .A(N565), .B(N564), .C(N636), .D(N569), .Y(N566) );
  NAND2X1TF U963 ( .A(N179), .B(N157), .Y(N587) );
  NOR4XLTF U964 ( .A(\RSHT_BITS[3] ), .B(N90), .C(N611), .D(N587), .Y(N568) );
  NAND2X1TF U965 ( .A(N576), .B(N586), .Y(N583) );
  NAND2X1TF U966 ( .A(N92), .B(N91), .Y(N585) );
  AOI2BB2X1TF U967 ( .B0(N593), .B1(N157), .A0N(N587), .A1N(N589), .Y(N581) );
  NAND4X1TF U968 ( .A(N94), .B(N631), .C(N630), .D(N629), .Y(N632) );
  NAND4X1TF U969 ( .A(N637), .B(N636), .C(N635), .D(N640), .Y(N697) );
  NAND3X1TF U970 ( .A(N752), .B(N648), .C(N647), .Y(N649) );
  AO22X1TF U971 ( .A0(DIVISION_REMA[4]), .A1(N731), .B0(N192), .B1(N786), .Y(
        N739) );
  AOI2BB1X1TF U972 ( .A0N(X_IN[1]), .A1N(N760), .B0(N759), .Y(N763) );
  NAND4X1TF U973 ( .A(N790), .B(N789), .C(N788), .D(N787), .Y(N791) );
  OAI221XLTF U974 ( .A0(\INDEX[2] ), .A1(N90), .B0(N124), .B1(\RSHT_BITS[3] ), 
        .C0(N813), .Y(N814) );
  OAI221XLTF U975 ( .A0(N129), .A1(N179), .B0(N156), .B1(N92), .C0(N815), .Y(
        N831) );
  NAND2X1TF U976 ( .A(N892), .B(N864), .Y(N861) );
  NAND2BX1TF U977 ( .AN(N816), .B(N861), .Y(N879) );
  NAND2X1TF U978 ( .A(N830), .B(N964), .Y(N865) );
  NAND3X1TF U979 ( .A(SIGN_Y), .B(N74), .C(N222), .Y(N838) );
  OAI2BB1X1TF U980 ( .A0N(N957), .A1N(N831), .B0(N830), .Y(N915) );
  NAND3X1TF U981 ( .A(N74), .B(N177), .C(N56), .Y(N972) );
  NAND4X1TF U982 ( .A(N222), .B(N177), .C(N56), .D(N962), .Y(N840) );
  NAND2X1TF U983 ( .A(N892), .B(N915), .Y(N940) );
  NAND3X1TF U984 ( .A(N904), .B(N903), .C(N902), .Y(N673) );
  NAND2X1TF U985 ( .A(N976), .B(N975), .Y(N668) );
  NAND2X1TF U986 ( .A(N979), .B(N978), .Y(N667) );
  NAND2X1TF U987 ( .A(SUM_AB[3]), .B(N83), .Y(N980) );
  NAND2X1TF U988 ( .A(N985), .B(N984), .Y(N665) );
  NAND2X1TF U989 ( .A(SUM_AB[5]), .B(N83), .Y(N986) );
  NAND2X1TF U990 ( .A(N991), .B(N990), .Y(N663) );
  NAND2X1TF U991 ( .A(SUM_AB[7]), .B(N83), .Y(N992) );
  NAND2X1TF U992 ( .A(N997), .B(N996), .Y(N661) );
  NAND2X1TF U993 ( .A(SUM_AB[9]), .B(N83), .Y(N998) );
  NAND2X1TF U994 ( .A(N1003), .B(N1002), .Y(N659) );
  NAND2X1TF U995 ( .A(SUM_AB[11]), .B(N83), .Y(N1004) );
endmodule


module SERIAL_CPU_8BIT_VG ( CLK, ENABLE, RST_N, START, I_DATAIN, D_DATAIN, 
        IS_I_ADDR, NXT, I_ADDR, D_ADDR, D_WE, D_DATAOUT, IO_STATUS, IO_CONTROL, 
        IO_DATAINA, IO_DATAINB, IO_DATAOUTA, IO_DATAOUTB, IO_OFFSET );
  input [7:0] I_DATAIN;
  input [7:0] D_DATAIN;
  output [1:0] NXT;
  output [8:0] I_ADDR;
  output [8:0] D_ADDR;
  output [7:0] D_DATAOUT;
  input [15:0] IO_STATUS;
  output [15:0] IO_CONTROL;
  input [15:0] IO_DATAINA;
  input [15:0] IO_DATAINB;
  output [15:0] IO_DATAOUTA;
  output [15:0] IO_DATAOUTB;
  output [15:0] IO_OFFSET;
  input CLK, ENABLE, RST_N, START;
  output IS_I_ADDR, D_WE;
  wire   \OPER1_R1[2] , \STATE[3] , N172, N173, N174, CF_BUF, N476, N477, N478,
         N479, N480, N481, N482, N483, N484, N485, N486, N487, N488, N489,
         N490, N491, N492, N510, N511, N512, N513, N514, N515, N516, N517,
         N518, N519, N520, N521, N522, N523, N524, N525, N594, N595, ZF, CF,
         N622, N402, N403, N404, N405, N406, N416, N418, N423, N435, N436,
         N437, N438, N439, N440, N441, N442, N443, N444, N445, N446, N447,
         N449, N450, N451, N453, N454, N455, N457, N458, N459, N461, N462,
         N463, N464, N466, N467, N468, N470, N471, N472, N474, N475, N4760,
         N4770, N4790, N4800, N4810, N4820, N4840, N4850, N4860, N4880, N4890,
         N4900, N4910, N493, N494, N495, N497, N498, N499, N500, N502, N503,
         N504, N505, N507, N508, N509, N5100, N5120, N5130, N5150, N5160,
         N5220, N5240, N5250, N526, N527, N528, N529, N530, N531, N532, N533,
         N534, N535, N536, N537, N538, N539, N557, N558, N559, N572, N574,
         N575, N598, N599, N600, N601, N602, N603, N604, N605, N606, N607,
         N608, N609, N610, N611, N612, N613, N616, N617, N618, N619, N620,
         N621, N6220, N623, N624, N625, N626, N627, N628, N629, N630, N631,
         N632, N633, N634, N635, N636, N637, N638, N639, N640, N641, N642,
         N643, N644, N645, N646, N647, N648, N649, N650, N651, N652, N653,
         N654, N655, N656, N657, N658, N659, N660, N661, N662, N663, N664,
         N665, N666, N667, N668, N669, N670, N671, N672, N673, N674, N675,
         N676, N677, N678, N679, N680, N681, N682, N683, N684, N685, N686,
         N687, N688, N689, N690, N691, N692, N693, N694, N695, N696, N808,
         N812, N813, N814, N815, N816, N864, N865, N927, N928, N929, N930,
         N931, N932, N933, N934, N935, N936, N937, N938, N939, N940, N941,
         N942, N943, N944, N945, N946, N947, N948, N949, N950, N951, N952,
         N953, N954, N955, N956, N957, N958, N959, N960, N961, N962, N963,
         N964, N965, N966, N967, N968, N969, N970, N971, N972, N973, N974,
         N975, N976, N977, N978, N979, N980, N981, N982, N983, N984, N985,
         N986, N987, N988, N989, N990, N991, N992, N993, N994, N995, N996,
         N997, N998, N999, N1000, N1001, N1002, N1003, N1004, N1005, N1006,
         N1007, N1008, SUB_X_292_4_N16, SUB_X_292_4_N15, SUB_X_292_4_N14,
         SUB_X_292_4_N13, SUB_X_292_4_N12, SUB_X_292_4_N11, SUB_X_292_4_N10,
         SUB_X_292_4_N9, SUB_X_292_4_N8, SUB_X_292_4_N7, SUB_X_292_4_N6,
         SUB_X_292_4_N5, SUB_X_292_4_N4, SUB_X_292_4_N3, SUB_X_292_4_N2,
         SUB_X_292_4_N1, ADD_X_292_3_N16, ADD_X_292_3_N15, ADD_X_292_3_N14,
         ADD_X_292_3_N13, ADD_X_292_3_N12, ADD_X_292_3_N11, ADD_X_292_3_N10,
         ADD_X_292_3_N9, ADD_X_292_3_N8, ADD_X_292_3_N7, ADD_X_292_3_N6,
         ADD_X_292_3_N5, ADD_X_292_3_N4, ADD_X_292_3_N3, ADD_X_292_3_N2, N1,
         N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N49, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166,
         N167, N168, N169, N170, N171, N1720, N1730, N1740, N175, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N190, N191, N192, N193, N194, N195, N196, N197, N198, N199,
         N200, N208, N209, N210, N211, N212, N213, N214, N215, N216, N217,
         N218, N219, N220, N221, N222, N223, N224, N225, N226, N227, N228,
         N229, N230, N231, N232, N233, N234, N235, N236, N237, N238, N239,
         N240, N241, N242, N243, N244, N245, N246, N247, N248, N249, N250,
         N251, N252, N253, N254, N255, N256, N257, N258, N259, N260, N261,
         N262, N263, N264, N265, N266, N267, N268, N269, N270, N271, N272,
         N273, N274, N275, N276, N277, N278, N279, N280, N281, N282, N283,
         N284, N285, N286, N287, N288, N289, N290, N291, N292, N293, N294,
         N295, N296, N297, N298, N299, N300, N301, N302, N303, N304, N305,
         N306, N307, N308, N309, N310, N311, N312, N313, N314, N315, N316,
         N317, N318, N319, N320, N321, N322, N323, N324, N325, N326, N327,
         N328, N329, N330, N331, N332, N333, N334, N335, N336, N337, N338,
         N339, N340, N341, N342, N343, N344, N345, N346, N347, N348, N349,
         N350, N351, N352, N353, N354, N355, N356, N357, N358, N359, N360,
         N361, N362, N363, N364, N365, N366, N367, N368, N369, N370, N371,
         N372, N373, N374, N375, N376, N377, N378, N379, N380, N381, N382,
         N383, N384, N385, N386, N387, N388, N389, N390, N391, N392, N393,
         N394, N395, N396, N397, N398, N399, N400, N401, N407, N408, N409,
         N410, N411, N412, N413, N414, N415, N417, N419, N420, N421, N422,
         N424, N425, N426, N427, N428, N429, N430, N431, N432, N433, N434,
         N448, N452, N456, N460, N465, N469, N473, N4780, N4830, N4870, N4920,
         N496, N501, N506, N5110, N5140, N5170, N5180, N5190, N5210, N5230,
         N540, N541, N542, N543, N544, N545, N546, N547, N548, N549, N550,
         N551, N552, N553, N554, N555, N556, N560, N561, N562, N563, N564,
         N565, N566, N567, N568, N569, N570, N571, N573, N576, N577, N578,
         N579, N580, N581, N582, N583, N584, N585, N586, N587, N588, N589,
         N590, N591, N592, N593, N5940, N5950, N596, N597, N614, N615, N697,
         N698, N699, N700, N701, N702, N703, N704, N705, N706, N707, N708,
         N709, N710, N711, N712, N713, N714, N715, N716, N717, N718, N719,
         N720, N721, N722, N723, N724, N725, N726, N727, N728, N729, N730,
         N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741,
         N742, N743, N744, N745, N746, N747, N748, N749, N750, N751, N752,
         N753, N754, N755, N756, N757, N758, N759, N760, N761, N762, N763,
         N764, N765, N766, N767, N768, N769, N770, N771, N772, N773, N774,
         N775, N776, N777, N778, N779, N780, N781, N782, N783, N784, N785,
         N786, N787, N788, N789, N790, N791, N792, N793, N794, N795, N796,
         N797, N798, N799, N800, N801, N802, N803, N804, N805, N806, N807,
         N809, N810, N811, N817, N818, N819, N820, N821, N822, N823, N824,
         N825, N826, N827, N828, N829, N830, N831, N832, N833, N834, N835,
         N836, N837, N838, N839, N840, N841, N842, N843, N844, N845, N846,
         N847, N848, N849, N850, N851, N852, N853, N854, N855, N856, N857,
         N858, N859, N860, N861, N862, N863, N866, N867, N868, N869, N870,
         N871, N872, N873, N874, N875, N876, N877, N878, N879, N880, N881,
         N882, N883, N884, N885, N886, N887, N888, N889, N890, N891, N892,
         N893, N894, N895, N896, N897, N898, N899, N900, N901, N902, N903,
         N904, N905, N906, N907, N908, N909, N910, N911, N912, N913, N914,
         N915, N916, N917, N918, N919, N920, N921, N922, N923, N924, N925,
         N926, N1009, N1010, N1011, N1012, N1013, N1014, N1015, N1016, N1017,
         N1018, N1019, N1020, N1021, N1022, N1023, N1024, N1025, N1026, N1027,
         N1028, N1029, N1030, N1031, N1032, N1033, N1034, N1035, N1036, N1037,
         N1038, N1039, N1040, N1041, N1042, N1043, N1044, N1045, N1046, N1047,
         N1048, N1049, N1050, N1051, N1052, N1053, N1054, N1055, N1056, N1057,
         N1058, N1059, N1060, N1061, N1062, N1063, N1064, N1065, N1066, N1067,
         N1068, N1069, N1070, N1071, N1072, N1073, N1074, N1075, N1076, N1077,
         N1078, N1079, N1080, N1081, N1082, N1083, N1084, N1085, N1086, N1087,
         N1088, N1089, N1090, N1091, N1092, N1093, N1094, N1095, N1096, N1097,
         N1098, N1099, N1100, N1101, N1102, N1103, N1104, N1105, N1106, N1107,
         N1108, N1109, N1110, N1111, N1112, N1113, N1114, N1115, N1116, N1117,
         N1118, N1119, N1120, N1121, N1122, N1123, N1124, N1125, N1126, N1127,
         N1128, N1129, N1130, N1131, N1132, N1133, N1134, N1135, N1136, N1137,
         N1138, N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1146, N1147,
         N1148, N1149, N1150, N1151, N1152, N1153, N1154, N1155, N1156, N1157,
         N1158, N1159, N1160, N1161, N1162, N1163, N1164, N1165, N1166, N1167,
         N1168, N1169, N1170, N1171, N1172, N1173, N1174, N1175, N1176, N1177,
         N1178, N1179, N1180, N1181, N1182, N1183, N1184, N1185, N1186, N1187,
         N1188, N1189, N1190, N1191, N1192, N1193, N1194, N1195, N1196, N1197,
         N1198;
  wire   [4:2] CODE_TYPE;
  wire   [2:0] OPER3_R3;
  wire   [3:0] NEXT_STATE;
  wire   [15:0] REG_A;
  wire   [15:0] REG_B;
  wire   [12:8] REG_C;

  DFFRX4TF \reg_A_reg[0]  ( .D(N499), .CK(CLK), .RN(RST_N), .Q(REG_A[0]), .QN(
        N222) );
  DFFRX4TF \reg_B_reg[0]  ( .D(N498), .CK(CLK), .RN(RST_N), .Q(REG_B[0]), .QN(
        N38) );
  CLKINVX6TF U551 ( .A(RST_N), .Y(N696) );
  DFFSX2TF \pc_reg[6]  ( .D(N808), .CK(CLK), .SN(RST_N), .Q(N245), .QN(
        I_ADDR[7]) );
  DFFSX2TF \pc_reg[4]  ( .D(N813), .CK(CLK), .SN(RST_N), .Q(N242), .QN(
        I_ADDR[5]) );
  DFFSX2TF \pc_reg[1]  ( .D(N816), .CK(CLK), .SN(RST_N), .Q(N241), .QN(
        I_ADDR[2]) );
  DFFSX2TF \pc_reg[0]  ( .D(N865), .CK(CLK), .SN(RST_N), .Q(N233), .QN(
        I_ADDR[1]) );
  DFFSX2TF \pc_reg[2]  ( .D(N815), .CK(CLK), .SN(RST_N), .Q(N216), .QN(
        I_ADDR[3]) );
  TLATXLTF cf_buf_reg ( .G(N594), .D(N595), .Q(CF_BUF) );
  TLATXLTF \nxt_reg[0]  ( .G(N172), .D(N173), .Q(NXT[0]) );
  TLATXLTF \nxt_reg[1]  ( .G(N172), .D(N174), .Q(NXT[1]) );
  DFFSX2TF \pc_reg[5]  ( .D(N812), .CK(CLK), .SN(RST_N), .QN(I_ADDR[6]) );
  DFFSX2TF \pc_reg[7]  ( .D(N864), .CK(CLK), .SN(RST_N), .QN(I_ADDR[8]) );
  DFFSX2TF \pc_reg[3]  ( .D(N814), .CK(CLK), .SN(RST_N), .QN(I_ADDR[4]) );
  DFFNSRX1TF \reg_C_reg[15]  ( .D(N497), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N416) );
  CMPR32X2TF \sub_x_292_4/U9  ( .A(N193), .B(REG_A[8]), .C(SUB_X_292_4_N9), 
        .CO(SUB_X_292_4_N8), .S(N518) );
  CMPR32X2TF \sub_x_292_4/U6  ( .A(N196), .B(REG_A[11]), .C(SUB_X_292_4_N6), 
        .CO(SUB_X_292_4_N5), .S(N521) );
  CMPR32X2TF \sub_x_292_4/U10  ( .A(N192), .B(REG_A[7]), .C(SUB_X_292_4_N10), 
        .CO(SUB_X_292_4_N9), .S(N517) );
  CMPR32X2TF \sub_x_292_4/U11  ( .A(N191), .B(REG_A[6]), .C(SUB_X_292_4_N11), 
        .CO(SUB_X_292_4_N10), .S(N516) );
  CMPR32X2TF \sub_x_292_4/U5  ( .A(N197), .B(REG_A[12]), .C(SUB_X_292_4_N5), 
        .CO(SUB_X_292_4_N4), .S(N522) );
  CMPR32X2TF \sub_x_292_4/U2  ( .A(N200), .B(REG_A[15]), .C(SUB_X_292_4_N2), 
        .CO(SUB_X_292_4_N1), .S(N525) );
  CMPR32X2TF \sub_x_292_4/U16  ( .A(N187), .B(REG_A[1]), .C(SUB_X_292_4_N16), 
        .CO(SUB_X_292_4_N15), .S(N511) );
  CMPR32X2TF \sub_x_292_4/U4  ( .A(N198), .B(REG_A[13]), .C(SUB_X_292_4_N4), 
        .CO(SUB_X_292_4_N3), .S(N523) );
  CMPR32X2TF \sub_x_292_4/U3  ( .A(N199), .B(REG_A[14]), .C(SUB_X_292_4_N3), 
        .CO(SUB_X_292_4_N2), .S(N524) );
  CMPR32X2TF \add_x_292_3/U5  ( .A(REG_A[12]), .B(REG_B[12]), .C(
        ADD_X_292_3_N5), .CO(ADD_X_292_3_N4), .S(N488) );
  CMPR32X2TF \add_x_292_3/U6  ( .A(REG_A[11]), .B(REG_B[11]), .C(
        ADD_X_292_3_N6), .CO(ADD_X_292_3_N5), .S(N487) );
  CMPR32X2TF \add_x_292_3/U7  ( .A(REG_A[10]), .B(REG_B[10]), .C(
        ADD_X_292_3_N7), .CO(ADD_X_292_3_N6), .S(N486) );
  CMPR32X2TF \add_x_292_3/U3  ( .A(REG_A[14]), .B(REG_B[14]), .C(
        ADD_X_292_3_N3), .CO(ADD_X_292_3_N2), .S(N490) );
  CMPR32X2TF \add_x_292_3/U16  ( .A(REG_A[1]), .B(REG_B[1]), .C(
        ADD_X_292_3_N16), .CO(ADD_X_292_3_N15), .S(N477) );
  CMPR32X2TF \add_x_292_3/U15  ( .A(REG_A[2]), .B(N135), .C(ADD_X_292_3_N15), 
        .CO(ADD_X_292_3_N14), .S(N478) );
  CMPR32X2TF \add_x_292_3/U14  ( .A(REG_A[3]), .B(REG_B[3]), .C(
        ADD_X_292_3_N14), .CO(ADD_X_292_3_N13), .S(N479) );
  CMPR32X2TF \add_x_292_3/U13  ( .A(REG_A[4]), .B(REG_B[4]), .C(
        ADD_X_292_3_N13), .CO(ADD_X_292_3_N12), .S(N480) );
  CMPR32X2TF \add_x_292_3/U12  ( .A(REG_A[5]), .B(REG_B[5]), .C(
        ADD_X_292_3_N12), .CO(ADD_X_292_3_N11), .S(N481) );
  CMPR32X2TF \add_x_292_3/U11  ( .A(REG_A[6]), .B(REG_B[6]), .C(
        ADD_X_292_3_N11), .CO(ADD_X_292_3_N10), .S(N482) );
  CMPR32X2TF \add_x_292_3/U10  ( .A(REG_A[7]), .B(REG_B[7]), .C(
        ADD_X_292_3_N10), .CO(ADD_X_292_3_N9), .S(N483) );
  CMPR32X2TF \add_x_292_3/U9  ( .A(REG_A[8]), .B(REG_B[8]), .C(ADD_X_292_3_N9), 
        .CO(ADD_X_292_3_N8), .S(N484) );
  CMPR32X2TF \add_x_292_3/U8  ( .A(REG_A[9]), .B(REG_B[9]), .C(ADD_X_292_3_N8), 
        .CO(ADD_X_292_3_N7), .S(N485) );
  CMPR32X2TF \add_x_292_3/U4  ( .A(REG_A[13]), .B(REG_B[13]), .C(
        ADD_X_292_3_N4), .CO(ADD_X_292_3_N3), .S(N489) );
  DFFNSRXLTF is_i_addr_reg ( .D(N1007), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        IS_I_ADDR), .QN(N250) );
  DFFNSRXLTF \reg_C_reg[13]  ( .D(N470), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N423) );
  DFFNSRXLTF \reg_C_reg[14]  ( .D(N4880), .CKN(CLK), .SN(1'b1), .RN(1'b1), 
        .QN(N418) );
  DFFNSRXLTF dw_reg ( .D(N622), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(D_WE) );
  DFFNSRXLTF \reg_C_reg[12]  ( .D(N507), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        REG_C[12]) );
  DFFNSRXLTF \reg_C_reg[11]  ( .D(N5120), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        REG_C[11]) );
  DFFNSRXLTF \reg_C_reg[9]  ( .D(N474), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        REG_C[9]) );
  DFFNSRXLTF \reg_C_reg[8]  ( .D(N461), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        REG_C[8]) );
  DFFNSRXLTF \reg_C_reg[10]  ( .D(N4790), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        REG_C[10]) );
  DFFRX2TF \reg_B_reg[1]  ( .D(N4890), .CK(CLK), .RN(RST_N), .Q(REG_B[1]), 
        .QN(N187) );
  DFFRX1TF \smdr_reg[8]  ( .D(N459), .CK(CLK), .RN(RST_N), .QN(N605) );
  DFFRX1TF \smdr_reg[6]  ( .D(N451), .CK(CLK), .RN(RST_N), .QN(N607) );
  DFFRX1TF \smdr_reg[4]  ( .D(N455), .CK(CLK), .RN(RST_N), .QN(N609) );
  DFFRX1TF \smdr_reg[3]  ( .D(N4820), .CK(CLK), .RN(RST_N), .QN(N610) );
  DFFRX1TF \smdr_reg[1]  ( .D(N4910), .CK(CLK), .RN(RST_N), .QN(N612) );
  DFFRX1TF \smdr_reg[0]  ( .D(N500), .CK(CLK), .RN(RST_N), .QN(N613) );
  DFFRX1TF \smdr_reg[5]  ( .D(N447), .CK(CLK), .RN(RST_N), .QN(N608) );
  DFFRX1TF \smdr_reg[15]  ( .D(N495), .CK(CLK), .RN(RST_N), .QN(N598) );
  DFFRX1TF \smdr_reg[14]  ( .D(N4860), .CK(CLK), .RN(RST_N), .QN(N599) );
  DFFRX1TF \smdr_reg[13]  ( .D(N468), .CK(CLK), .RN(RST_N), .QN(N600) );
  DFFRX1TF \smdr_reg[12]  ( .D(N505), .CK(CLK), .RN(RST_N), .QN(N601) );
  DFFRX1TF \smdr_reg[11]  ( .D(N5100), .CK(CLK), .RN(RST_N), .QN(N602) );
  DFFRX1TF \smdr_reg[10]  ( .D(N4770), .CK(CLK), .RN(RST_N), .QN(N603) );
  DFFRX1TF \smdr_reg[9]  ( .D(N472), .CK(CLK), .RN(RST_N), .QN(N604) );
  DFFRX1TF \smdr_reg[7]  ( .D(N435), .CK(CLK), .RN(RST_N), .QN(N606) );
  DFFRX1TF \smdr_reg[2]  ( .D(N464), .CK(CLK), .RN(RST_N), .QN(N611) );
  DFFRX1TF nf_reg ( .D(N437), .CK(CLK), .RN(RST_N), .QN(N244) );
  DFFRX1TF \id_ir_reg[7]  ( .D(N532), .CK(CLK), .RN(RST_N), .QN(N406) );
  DFFRX1TF \id_ir_reg[3]  ( .D(N536), .CK(CLK), .RN(RST_N), .QN(N402) );
  DFFRX1TF \id_ir_reg[6]  ( .D(N533), .CK(CLK), .RN(RST_N), .QN(N405) );
  DFFRX1TF \id_ir_reg[5]  ( .D(N534), .CK(CLK), .RN(RST_N), .QN(N404) );
  DFFRX1TF \gr_reg[0][15]  ( .D(N958), .CK(CLK), .RN(RST_N), .QN(N680) );
  DFFRX1TF \gr_reg[0][14]  ( .D(N959), .CK(CLK), .RN(RST_N), .QN(N681) );
  DFFRX1TF \gr_reg[0][13]  ( .D(N960), .CK(CLK), .RN(RST_N), .QN(N682) );
  DFFRX1TF \gr_reg[4][15]  ( .D(N1006), .CK(CLK), .RN(RST_N), .QN(N616) );
  DFFRX1TF \gr_reg[4][14]  ( .D(N927), .CK(CLK), .RN(RST_N), .QN(N617) );
  DFFRX1TF \gr_reg[4][13]  ( .D(N928), .CK(CLK), .RN(RST_N), .QN(N618) );
  DFFRX1TF \gr_reg[2][15]  ( .D(N942), .CK(CLK), .RN(RST_N), .QN(N648) );
  DFFRX1TF \gr_reg[2][14]  ( .D(N943), .CK(CLK), .RN(RST_N), .QN(N649) );
  DFFRX1TF \gr_reg[2][13]  ( .D(N944), .CK(CLK), .RN(RST_N), .QN(N650) );
  DFFRX1TF \gr_reg[1][15]  ( .D(N950), .CK(CLK), .RN(RST_N), .QN(N664) );
  DFFRX1TF \gr_reg[1][14]  ( .D(N951), .CK(CLK), .RN(RST_N), .QN(N665) );
  DFFRX1TF \gr_reg[1][13]  ( .D(N952), .CK(CLK), .RN(RST_N), .QN(N666) );
  DFFRX1TF \gr_reg[0][12]  ( .D(N961), .CK(CLK), .RN(RST_N), .QN(N683) );
  DFFRX1TF \gr_reg[0][11]  ( .D(N962), .CK(CLK), .RN(RST_N), .QN(N684) );
  DFFRX1TF \gr_reg[0][10]  ( .D(N963), .CK(CLK), .RN(RST_N), .QN(N685) );
  DFFRX1TF \gr_reg[0][9]  ( .D(N964), .CK(CLK), .RN(RST_N), .QN(N686) );
  DFFRX1TF \gr_reg[0][8]  ( .D(N965), .CK(CLK), .RN(RST_N), .QN(N687) );
  DFFRX1TF \gr_reg[0][4]  ( .D(N1001), .CK(CLK), .RN(RST_N), .QN(N691) );
  DFFRX1TF \gr_reg[0][3]  ( .D(N1002), .CK(CLK), .RN(RST_N), .QN(N692) );
  DFFRX1TF \gr_reg[0][2]  ( .D(N1003), .CK(CLK), .RN(RST_N), .QN(N693) );
  DFFRX1TF \gr_reg[0][1]  ( .D(N1004), .CK(CLK), .RN(RST_N), .QN(N694) );
  DFFRX1TF \gr_reg[0][0]  ( .D(N1005), .CK(CLK), .RN(RST_N), .QN(N695) );
  DFFRX1TF \gr_reg[4][12]  ( .D(N929), .CK(CLK), .RN(RST_N), .QN(N619) );
  DFFRX1TF \gr_reg[4][11]  ( .D(N930), .CK(CLK), .RN(RST_N), .QN(N620) );
  DFFRX1TF \gr_reg[4][10]  ( .D(N931), .CK(CLK), .RN(RST_N), .QN(N621) );
  DFFRX1TF \gr_reg[0][7]  ( .D(N998), .CK(CLK), .RN(RST_N), .QN(N688) );
  DFFRX1TF \gr_reg[0][6]  ( .D(N999), .CK(CLK), .RN(RST_N), .QN(N689) );
  DFFRX1TF \gr_reg[0][5]  ( .D(N1000), .CK(CLK), .RN(RST_N), .QN(N690) );
  DFFRX1TF \gr_reg[1][12]  ( .D(N953), .CK(CLK), .RN(RST_N), .QN(N667) );
  DFFRX1TF \gr_reg[1][11]  ( .D(N954), .CK(CLK), .RN(RST_N), .QN(N668) );
  DFFRX1TF \gr_reg[1][10]  ( .D(N955), .CK(CLK), .RN(RST_N), .QN(N669) );
  DFFRX1TF \gr_reg[1][9]  ( .D(N956), .CK(CLK), .RN(RST_N), .QN(N670) );
  DFFRX1TF \gr_reg[1][8]  ( .D(N957), .CK(CLK), .RN(RST_N), .QN(N671) );
  DFFRX1TF \gr_reg[1][7]  ( .D(N990), .CK(CLK), .RN(RST_N), .QN(N672) );
  DFFRX1TF cf_reg ( .D(N5220), .CK(CLK), .RN(RST_N), .Q(CF) );
  DFFRX1TF \reg_B_reg[2]  ( .D(N462), .CK(CLK), .RN(RST_N), .Q(N40), .QN(N134)
         );
  DFFRX2TF \state_reg[3]  ( .D(NEXT_STATE[3]), .CK(CLK), .RN(RST_N), .Q(
        \STATE[3] ), .QN(N232) );
  DFFRX2TF \state_reg[0]  ( .D(NEXT_STATE[0]), .CK(CLK), .RN(RST_N), .Q(N215), 
        .QN(N559) );
  DFFRX2TF \state_reg[2]  ( .D(NEXT_STATE[2]), .CK(CLK), .RN(RST_N), .Q(N221), 
        .QN(N557) );
  DFFRX2TF \state_reg[1]  ( .D(NEXT_STATE[1]), .CK(CLK), .RN(RST_N), .Q(N211), 
        .QN(N558) );
  DFFRX2TF \reg_A_reg[4]  ( .D(N454), .CK(CLK), .RN(RST_N), .Q(REG_A[4]), .QN(
        N237) );
  DFFRX2TF \reg_B_reg[13]  ( .D(N441), .CK(CLK), .RN(RST_N), .Q(REG_B[13]), 
        .QN(N198) );
  DFFRX2TF \reg_A_reg[14]  ( .D(N4850), .CK(CLK), .RN(RST_N), .Q(REG_A[14]), 
        .QN(N210) );
  DFFRX2TF \reg_A_reg[9]  ( .D(N471), .CK(CLK), .RN(RST_N), .Q(REG_A[9]), .QN(
        N220) );
  DFFRX2TF \reg_A_reg[7]  ( .D(N5130), .CK(CLK), .RN(RST_N), .Q(REG_A[7]), 
        .QN(N224) );
  DFFRX2TF \reg_A_reg[3]  ( .D(N4810), .CK(CLK), .RN(RST_N), .Q(REG_A[3]), 
        .QN(N219) );
  DFFRX2TF \reg_A_reg[15]  ( .D(N494), .CK(CLK), .RN(RST_N), .Q(REG_A[15]), 
        .QN(N229) );
  DFFRX2TF \reg_A_reg[13]  ( .D(N467), .CK(CLK), .RN(RST_N), .Q(REG_A[13]), 
        .QN(N226) );
  DFFRX2TF \reg_A_reg[12]  ( .D(N504), .CK(CLK), .RN(RST_N), .Q(REG_A[12]), 
        .QN(N227) );
  DFFRX2TF \reg_A_reg[11]  ( .D(N509), .CK(CLK), .RN(RST_N), .Q(REG_A[11]), 
        .QN(N231) );
  DFFRX2TF \reg_A_reg[10]  ( .D(N4760), .CK(CLK), .RN(RST_N), .Q(REG_A[10]), 
        .QN(N223) );
  DFFRX2TF \reg_A_reg[8]  ( .D(N458), .CK(CLK), .RN(RST_N), .Q(REG_A[8]), .QN(
        N239) );
  DFFRX2TF \reg_A_reg[2]  ( .D(N463), .CK(CLK), .RN(RST_N), .Q(REG_A[2]), .QN(
        N225) );
  DFFRX2TF \reg_A_reg[1]  ( .D(N4900), .CK(CLK), .RN(RST_N), .Q(REG_A[1]), 
        .QN(N208) );
  DFFRX2TF \reg_A_reg[6]  ( .D(N450), .CK(CLK), .RN(RST_N), .Q(REG_A[6]), .QN(
        N240) );
  DFFRX2TF \reg_A_reg[5]  ( .D(N446), .CK(CLK), .RN(RST_N), .Q(REG_A[5]), .QN(
        N209) );
  DFFRX2TF \reg_B_reg[15]  ( .D(N438), .CK(CLK), .RN(RST_N), .Q(REG_B[15]), 
        .QN(N200) );
  DFFRX2TF \reg_B_reg[14]  ( .D(N439), .CK(CLK), .RN(RST_N), .Q(REG_B[14]), 
        .QN(N199) );
  DFFRX2TF \reg_B_reg[8]  ( .D(N442), .CK(CLK), .RN(RST_N), .Q(REG_B[8]), .QN(
        N193) );
  DFFRX2TF \reg_B_reg[4]  ( .D(N443), .CK(CLK), .RN(RST_N), .Q(REG_B[4]), .QN(
        N189) );
  DFFRX2TF \reg_B_reg[7]  ( .D(N5160), .CK(CLK), .RN(RST_N), .Q(REG_B[7]), 
        .QN(N192) );
  DFFRX2TF \reg_B_reg[6]  ( .D(N444), .CK(CLK), .RN(RST_N), .Q(REG_B[6]), .QN(
        N191) );
  DFFRX2TF \reg_B_reg[5]  ( .D(N445), .CK(CLK), .RN(RST_N), .Q(REG_B[5]), .QN(
        N190) );
  DFFRX2TF \reg_B_reg[3]  ( .D(N4800), .CK(CLK), .RN(RST_N), .Q(REG_B[3]), 
        .QN(N188) );
  DFFRX2TF \reg_B_reg[12]  ( .D(N503), .CK(CLK), .RN(RST_N), .Q(REG_B[12]), 
        .QN(N197) );
  DFFRX2TF \reg_B_reg[11]  ( .D(N508), .CK(CLK), .RN(RST_N), .Q(REG_B[11]), 
        .QN(N196) );
  DFFRX2TF \reg_B_reg[10]  ( .D(N475), .CK(CLK), .RN(RST_N), .Q(REG_B[10]), 
        .QN(N195) );
  DFFRX2TF \reg_B_reg[9]  ( .D(N440), .CK(CLK), .RN(RST_N), .Q(REG_B[9]), .QN(
        N194) );
  DFFRX2TF zf_reg ( .D(N436), .CK(CLK), .RN(RST_N), .Q(ZF), .QN(N246) );
  DFFRX2TF \id_ir_reg[4]  ( .D(N535), .CK(CLK), .RN(RST_N), .Q(N236), .QN(N403) );
  DFFRX2TF \id_ir_reg[15]  ( .D(N5240), .CK(CLK), .RN(RST_N), .Q(CODE_TYPE[4]), 
        .QN(N212) );
  DFFRX2TF \id_ir_reg[11]  ( .D(N528), .CK(CLK), .RN(RST_N), .Q(N218), .QN(
        N572) );
  DFFRX2TF \id_ir_reg[2]  ( .D(N537), .CK(CLK), .RN(RST_N), .Q(OPER3_R3[2]), 
        .QN(N213) );
  DFFRX2TF \id_ir_reg[1]  ( .D(N538), .CK(CLK), .RN(RST_N), .Q(OPER3_R3[1]), 
        .QN(N217) );
  DFFRX2TF \id_ir_reg[0]  ( .D(N539), .CK(CLK), .RN(RST_N), .Q(OPER3_R3[0]), 
        .QN(N235) );
  DFFRX2TF \id_ir_reg[14]  ( .D(N5250), .CK(CLK), .RN(RST_N), .Q(CODE_TYPE[3]), 
        .QN(N228) );
  DFFRX2TF \id_ir_reg[13]  ( .D(N526), .CK(CLK), .RN(RST_N), .Q(CODE_TYPE[2]), 
        .QN(N214) );
  DFFRX2TF \id_ir_reg[10]  ( .D(N529), .CK(CLK), .RN(RST_N), .Q(\OPER1_R1[2] ), 
        .QN(N234) );
  DFFRX2TF \id_ir_reg[8]  ( .D(N531), .CK(CLK), .RN(RST_N), .Q(N243), .QN(N575) );
  DFFRX2TF \gr_reg[3][15]  ( .D(N934), .CK(CLK), .RN(RST_N), .Q(N249), .QN(
        N632) );
  DFFRX2TF \gr_reg[3][14]  ( .D(N935), .CK(CLK), .RN(RST_N), .Q(N248), .QN(
        N633) );
  DFFRX2TF \gr_reg[3][13]  ( .D(N936), .CK(CLK), .RN(RST_N), .Q(N247), .QN(
        N634) );
  DFFRX2TF \gr_reg[4][9]  ( .D(N932), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[9]), 
        .QN(N6220) );
  DFFRX2TF \gr_reg[4][8]  ( .D(N933), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[8]), 
        .QN(N623) );
  DFFRX2TF \gr_reg[4][4]  ( .D(N969), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[4]), 
        .QN(N627) );
  DFFRX2TF \gr_reg[4][3]  ( .D(N970), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[3]), 
        .QN(N628) );
  DFFRX2TF \gr_reg[4][2]  ( .D(N971), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[2]), 
        .QN(N629) );
  DFFRX2TF \gr_reg[4][1]  ( .D(N972), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[1]), 
        .QN(N630) );
  DFFRX2TF \gr_reg[4][0]  ( .D(N973), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[0]), 
        .QN(N631) );
  DFFRX2TF \gr_reg[4][7]  ( .D(N966), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[7]), 
        .QN(N624) );
  DFFRX2TF \gr_reg[4][6]  ( .D(N967), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[6]), 
        .QN(N625) );
  DFFRX2TF \gr_reg[4][5]  ( .D(N968), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[5]), 
        .QN(N626) );
  DFFRX2TF \gr_reg[3][12]  ( .D(N937), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTB[12]), .QN(N635) );
  DFFRX2TF \gr_reg[3][11]  ( .D(N938), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTB[11]), .QN(N636) );
  DFFRX2TF \gr_reg[3][10]  ( .D(N939), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTB[10]), .QN(N637) );
  DFFRX2TF \gr_reg[3][9]  ( .D(N940), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[9]), 
        .QN(N638) );
  DFFRX2TF \gr_reg[3][8]  ( .D(N941), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[8]), 
        .QN(N639) );
  DFFRX2TF \gr_reg[2][12]  ( .D(N945), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTA[12]), .QN(N651) );
  DFFRX2TF \gr_reg[2][11]  ( .D(N946), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTA[11]), .QN(N652) );
  DFFRX2TF \gr_reg[2][10]  ( .D(N947), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTA[10]), .QN(N653) );
  DFFRX2TF \gr_reg[2][9]  ( .D(N948), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[9]), 
        .QN(N654) );
  DFFRX2TF \gr_reg[2][8]  ( .D(N949), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[8]), 
        .QN(N655) );
  DFFRX2TF \gr_reg[3][4]  ( .D(N977), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[4]), 
        .QN(N643) );
  DFFRX2TF \gr_reg[3][3]  ( .D(N978), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[3]), 
        .QN(N644) );
  DFFRX2TF \gr_reg[3][2]  ( .D(N979), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[2]), 
        .QN(N645) );
  DFFRX2TF \gr_reg[3][1]  ( .D(N980), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[1]), 
        .QN(N646) );
  DFFRX2TF \gr_reg[3][0]  ( .D(N981), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[0]), 
        .QN(N647) );
  DFFRX2TF \gr_reg[2][4]  ( .D(N985), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[4]), 
        .QN(N659) );
  DFFRX2TF \gr_reg[2][3]  ( .D(N986), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[3]), 
        .QN(N660) );
  DFFRX2TF \gr_reg[2][2]  ( .D(N987), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[2]), 
        .QN(N661) );
  DFFRX2TF \gr_reg[2][1]  ( .D(N988), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[1]), 
        .QN(N662) );
  DFFRX2TF \gr_reg[2][0]  ( .D(N989), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[0]), 
        .QN(N663) );
  DFFRX2TF \gr_reg[3][7]  ( .D(N974), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[7]), 
        .QN(N640) );
  DFFRX2TF \gr_reg[3][6]  ( .D(N975), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[6]), 
        .QN(N641) );
  DFFRX2TF \gr_reg[3][5]  ( .D(N976), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[5]), 
        .QN(N642) );
  DFFRX2TF \gr_reg[2][7]  ( .D(N982), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[7]), 
        .QN(N656) );
  DFFRX2TF \gr_reg[2][6]  ( .D(N983), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[6]), 
        .QN(N657) );
  DFFRX2TF \gr_reg[2][5]  ( .D(N984), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[5]), 
        .QN(N658) );
  DFFRX2TF \gr_reg[1][4]  ( .D(N993), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[4]), 
        .QN(N675) );
  DFFRX2TF \gr_reg[1][3]  ( .D(N994), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[3]), 
        .QN(N676) );
  DFFRX2TF \gr_reg[1][2]  ( .D(N995), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[2]), 
        .QN(N677) );
  DFFRX2TF \gr_reg[1][1]  ( .D(N996), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[1]), 
        .QN(N678) );
  DFFRX2TF \gr_reg[1][0]  ( .D(N997), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[0]), 
        .QN(N679) );
  DFFRX2TF \gr_reg[1][6]  ( .D(N991), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[6]), 
        .QN(N673) );
  DFFRX2TF \gr_reg[1][5]  ( .D(N992), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[5]), 
        .QN(N674) );
  DFFNSRX2TF lowest_bit_reg ( .D(N1008), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        I_ADDR[0]), .QN(N230) );
  DFFRX2TF \id_ir_reg[9]  ( .D(N530), .CK(CLK), .RN(RST_N), .Q(N747), .QN(N574) );
  DFFNSRX2TF \reg_C_reg[2]  ( .D(N466), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[3]) );
  DFFNSRX2TF \reg_C_reg[4]  ( .D(N457), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[5]) );
  DFFNSRX2TF \reg_C_reg[6]  ( .D(N453), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[7]) );
  DFFNSRX2TF \reg_C_reg[5]  ( .D(N449), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[6]) );
  DFFNSRX2TF \reg_C_reg[1]  ( .D(N493), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[2]) );
  DFFNSRX2TF \reg_C_reg[3]  ( .D(N4840), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[4]) );
  DFFNSRX1TF \reg_C_reg[0]  ( .D(N502), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[1]) );
  DFFNSRX2TF \reg_C_reg[7]  ( .D(N5150), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[8]) );
  DFFRX2TF \id_ir_reg[12]  ( .D(N527), .CK(CLK), .RN(RST_N), .Q(N258), .QN(N39) );
  NAND2X1TF U3 ( .A(N420), .B(N188), .Y(N342) );
  OAI21X1TF U4 ( .A0(N396), .A1(N140), .B0(N395), .Y(N502) );
  XOR2X1TF U5 ( .A(N391), .B(N390), .Y(N396) );
  OAI21X1TF U6 ( .A0(N138), .A1(N237), .B0(N841), .Y(N1) );
  NOR3X1TF U7 ( .A(N839), .B(N840), .C(N1), .Y(N860) );
  NOR3BX1TF U8 ( .AN(N743), .B(N559), .C(\STATE[3] ), .Y(N421) );
  AO21X1TF U9 ( .A0(N259), .A1(N196), .B0(N136), .Y(N2) );
  AOI22X1TF U10 ( .A0(REG_A[11]), .A1(N424), .B0(N260), .B1(N231), .Y(N3) );
  AOI21X1TF U11 ( .A0(N149), .A1(N3), .B0(N196), .Y(N4) );
  AOI2BB2X1TF U12 ( .B0(N351), .B1(N771), .A0N(N820), .A1N(N848), .Y(N5) );
  OA22X1TF U13 ( .A0(N845), .A1(N810), .B0(N806), .B1(N885), .Y(N6) );
  OAI211X1TF U14 ( .A0(N772), .A1(N878), .B0(N5), .C0(N6), .Y(N7) );
  AOI211X1TF U15 ( .A0(REG_A[11]), .A1(N2), .B0(N4), .C0(N7), .Y(N8) );
  OAI2BB1X1TF U16 ( .A0N(N521), .A1N(N252), .B0(N8), .Y(N9) );
  AOI21X1TF U17 ( .A0(N253), .A1(N487), .B0(N9), .Y(N398) );
  NAND2BX1TF U18 ( .AN(N891), .B(N1014), .Y(N10) );
  OAI211X1TF U19 ( .A0(N1016), .A1(N426), .B0(N1015), .C0(N10), .Y(N1026) );
  NOR4XLTF U20 ( .A(N1195), .B(N370), .C(N371), .D(N376), .Y(N11) );
  NAND4X1TF U21 ( .A(N11), .B(N400), .C(N410), .D(N412), .Y(N12) );
  NOR4XLTF U22 ( .A(N383), .B(N407), .C(N378), .D(N12), .Y(N13) );
  AND4X1TF U23 ( .A(N13), .B(N387), .C(N397), .D(N398), .Y(N14) );
  NAND4X1TF U24 ( .A(N14), .B(N417), .C(N419), .D(N415), .Y(N15) );
  OAI2BB2XLTF U25 ( .B0(N391), .B1(N15), .A0N(N1195), .A1N(ZF), .Y(N436) );
  OAI222X1TF U26 ( .A0(N807), .A1(N848), .B0(N806), .B1(N878), .C0(N810), .C1(
        N851), .Y(N16) );
  AOI32X1TF U27 ( .A0(N422), .A1(REG_A[7]), .A2(N192), .B0(N136), .B1(REG_A[7]), .Y(N17) );
  OAI21X1TF U28 ( .A0(N820), .A1(N845), .B0(N17), .Y(N18) );
  AOI211X1TF U29 ( .A0(N339), .A1(N351), .B0(N16), .C0(N18), .Y(N19) );
  AOI22X1TF U30 ( .A0(REG_A[7]), .A1(N168), .B0(N260), .B1(N224), .Y(N20) );
  AOI32X1TF U31 ( .A0(N149), .A1(N19), .A2(N20), .B0(N192), .B1(N19), .Y(N21)
         );
  AO21X1TF U32 ( .A0(N517), .A1(N252), .B0(N21), .Y(N22) );
  AOI21X1TF U33 ( .A0(N363), .A1(N483), .B0(N22), .Y(N400) );
  OAI22X1TF U34 ( .A0(N680), .A1(N1184), .B0(N1160), .B1(N406), .Y(N23) );
  OAI22XLTF U35 ( .A0(N185), .A1(N632), .B0(N664), .B1(N1186), .Y(N24) );
  OAI22XLTF U36 ( .A0(N616), .A1(N159), .B0(N648), .B1(N1189), .Y(N25) );
  NOR3X1TF U37 ( .A(N23), .B(N24), .C(N25), .Y(N26) );
  OAI21X1TF U38 ( .A0(N200), .A1(N49), .B0(N26), .Y(N438) );
  AOI2BB2X1TF U39 ( .B0(N1182), .B1(IO_DATAINA[10]), .A0N(N387), .A1N(N139), 
        .Y(N27) );
  AOI22X1TF U40 ( .A0(REG_C[10]), .A1(N1180), .B0(IO_DATAINB[10]), .B1(N409), 
        .Y(N28) );
  OAI211X1TF U41 ( .A0(N397), .A1(N142), .B0(N27), .C0(N28), .Y(N4790) );
  AOI2BB2X1TF U42 ( .B0(N1182), .B1(IO_DATAINA[11]), .A0N(N397), .A1N(N139), 
        .Y(N29) );
  AOI22X1TF U43 ( .A0(REG_C[11]), .A1(N1180), .B0(IO_DATAINB[11]), .B1(N254), 
        .Y(N30) );
  OAI211X1TF U44 ( .A0(N398), .A1(N142), .B0(N29), .C0(N30), .Y(N5120) );
  OA21XLTF U45 ( .A0(N716), .A1(I_ADDR[4]), .B0(N717), .Y(N31) );
  AOI222XLTF U46 ( .A0(I_ADDR[4]), .A1(N722), .B0(N729), .B1(D_ADDR[4]), .C0(
        N720), .C1(N31), .Y(N814) );
  AOI2BB1X1TF U47 ( .A0N(N138), .A1N(N848), .B0(N5140), .Y(N327) );
  OAI21X1TF U48 ( .A0(N785), .A1(N220), .B0(N756), .Y(N32) );
  NOR3X1TF U49 ( .A(N754), .B(N755), .C(N32), .Y(N790) );
  AOI2BB2X1TF U50 ( .B0(N236), .B1(N1031), .A0N(N1035), .A1N(N1030), .Y(N156)
         );
  AOI2BB2X1TF U51 ( .B0(N1182), .B1(IO_DATAINA[12]), .A0N(N398), .A1N(N139), 
        .Y(N33) );
  AOI22X1TF U52 ( .A0(REG_C[12]), .A1(N1180), .B0(IO_DATAINB[12]), .B1(N254), 
        .Y(N34) );
  OAI211X1TF U53 ( .A0(N417), .A1(N142), .B0(N33), .C0(N34), .Y(N507) );
  OA21XLTF U54 ( .A0(N721), .A1(I_ADDR[6]), .B0(N726), .Y(N35) );
  AOI222XLTF U55 ( .A0(I_ADDR[6]), .A1(N722), .B0(N729), .B1(D_ADDR[6]), .C0(
        N720), .C1(N35), .Y(N812) );
  CLKINVX1TF U56 ( .A(N252), .Y(N36) );
  OAI22X1TF U57 ( .A0(SUB_X_292_4_N1), .A1(N36), .B0(N37), .B1(N542), .Y(N595)
         );
  CLKINVX1TF U58 ( .A(N492), .Y(N37) );
  OR3X1TF U59 ( .A(N1016), .B(N892), .C(N151), .Y(N883) );
  CLKBUFX2TF U60 ( .A(N1188), .Y(N49) );
  INVX1TF U79 ( .A(N860), .Y(N868) );
  CLKINVX4TF U80 ( .A(N422), .Y(N132) );
  OR3X1TF U81 ( .A(N752), .B(N890), .C(N746), .Y(N1168) );
  CLKINVX2TF U82 ( .A(N562), .Y(N271) );
  NAND2XLTF U83 ( .A(N426), .B(CODE_TYPE[3]), .Y(N893) );
  INVX2TF U84 ( .A(N258), .Y(N151) );
  AO22X1TF U85 ( .A0(N1033), .A1(N1032), .B0(N403), .B1(N1031), .Y(N1175) );
  OAI22X1TF U86 ( .A0(N234), .A1(N1035), .B0(N1034), .B1(N405), .Y(N1174) );
  OR2X2TF U87 ( .A(N1027), .B(N541), .Y(N858) );
  INVX2TF U88 ( .A(N900), .Y(N901) );
  OAI211XLTF U89 ( .A0(N1044), .A1(N1016), .B0(N560), .C0(N556), .Y(N561) );
  CLKINVX1TF U90 ( .A(N734), .Y(N735) );
  NAND2XLTF U91 ( .A(N427), .B(REG_A[5]), .Y(N774) );
  INVX2TF U92 ( .A(N137), .Y(N427) );
  ADDFHX2TF U93 ( .A(N133), .B(REG_A[2]), .CI(SUB_X_292_4_N15), .CO(
        SUB_X_292_4_N14), .S(N512) );
  INVX4TF U94 ( .A(N135), .Y(N133) );
  CMPR22X2TF U95 ( .A(REG_B[0]), .B(REG_A[0]), .CO(ADD_X_292_3_N16), .S(N476)
         );
  OAI222X1TF U96 ( .A0(N142), .A1(N388), .B0(N140), .B1(N415), .C0(N416), .C1(
        N251), .Y(N497) );
  XOR2X2TF U97 ( .A(N419), .B(N389), .Y(N390) );
  OA22X1TF U98 ( .A0(N412), .A1(N140), .B0(N413), .B1(N142), .Y(N1129) );
  AOI22X1TF U99 ( .A0(N701), .A1(N702), .B0(N639), .B1(N699), .Y(N941) );
  AOI22X1TF U100 ( .A0(N701), .A1(N706), .B0(N635), .B1(N699), .Y(N937) );
  AOI22X1TF U101 ( .A0(N701), .A1(N704), .B0(N637), .B1(N699), .Y(N939) );
  AOI22X1TF U102 ( .A0(N701), .A1(N705), .B0(N636), .B1(N699), .Y(N938) );
  AOI22X1TF U103 ( .A0(N697), .A1(N702), .B0(N655), .B1(N615), .Y(N949) );
  AOI22X1TF U104 ( .A0(N614), .A1(N706), .B0(N667), .B1(N597), .Y(N953) );
  AOI22X1TF U105 ( .A0(N697), .A1(N704), .B0(N653), .B1(N615), .Y(N947) );
  AOI22X1TF U106 ( .A0(N573), .A1(N588), .B0(N656), .B1(N571), .Y(N982) );
  AOI22X1TF U107 ( .A0(N573), .A1(N581), .B0(N662), .B1(N571), .Y(N988) );
  AOI22X1TF U108 ( .A0(N697), .A1(N706), .B0(N651), .B1(N615), .Y(N945) );
  AOI22X1TF U109 ( .A0(N614), .A1(N702), .B0(N671), .B1(N597), .Y(N957) );
  AOI22X1TF U110 ( .A0(N573), .A1(N585), .B0(N658), .B1(N571), .Y(N984) );
  AOI22X1TF U111 ( .A0(N697), .A1(N705), .B0(N652), .B1(N615), .Y(N946) );
  AOI22X1TF U112 ( .A0(N614), .A1(N704), .B0(N669), .B1(N597), .Y(N955) );
  NOR4XLTF U113 ( .A(N834), .B(N359), .C(N835), .D(N358), .Y(N360) );
  OAI22X1TF U114 ( .A0(N682), .A1(N184), .B0(N650), .B1(N181), .Y(N1081) );
  OAI22X1TF U115 ( .A0(N686), .A1(N184), .B0(N654), .B1(N181), .Y(N1087) );
  OAI22X1TF U116 ( .A0(N163), .A1(N605), .B0(N671), .B1(N177), .Y(N1064) );
  OAI22X1TF U117 ( .A0(N687), .A1(N183), .B0(N655), .B1(N180), .Y(N1063) );
  NAND3XLTF U118 ( .A(N543), .B(N859), .C(N542), .Y(N594) );
  OAI22X1TF U119 ( .A0(N695), .A1(N183), .B0(N663), .B1(N180), .Y(N1146) );
  OAI22X1TF U120 ( .A0(N693), .A1(N184), .B0(N661), .B1(N181), .Y(N1073) );
  OAI22X1TF U121 ( .A0(N161), .A1(N607), .B0(N673), .B1(N177), .Y(N1051) );
  OAI22X1TF U122 ( .A0(N685), .A1(N184), .B0(N653), .B1(N181), .Y(N1097) );
  OAI22X1TF U123 ( .A0(N688), .A1(N183), .B0(N656), .B1(N180), .Y(N748) );
  OAI22X1TF U124 ( .A0(N162), .A1(N609), .B0(N675), .B1(N177), .Y(N1057) );
  OAI22X1TF U125 ( .A0(N681), .A1(N184), .B0(N649), .B1(N181), .Y(N1115) );
  OAI22X1TF U126 ( .A0(N684), .A1(N184), .B0(N652), .B1(N181), .Y(N1169) );
  OAI22X1TF U127 ( .A0(N691), .A1(N183), .B0(N659), .B1(N180), .Y(N1056) );
  OAI22X1TF U128 ( .A0(N163), .A1(N613), .B0(N679), .B1(N177), .Y(N1147) );
  OAI22X1TF U129 ( .A0(N692), .A1(N183), .B0(N660), .B1(N180), .Y(N1107) );
  OAI22X1TF U130 ( .A0(N683), .A1(N184), .B0(N651), .B1(N181), .Y(N1157) );
  OAI22X1TF U131 ( .A0(N638), .A1(N1187), .B0(N670), .B1(N1186), .Y(N908) );
  AO22X1TF U132 ( .A0(N236), .A1(N1029), .B0(N1028), .B1(N1032), .Y(N1173) );
  OAI22X1TF U133 ( .A0(N689), .A1(N183), .B0(N657), .B1(N180), .Y(N1050) );
  OAI22X1TF U134 ( .A0(N162), .A1(N610), .B0(N676), .B1(N177), .Y(N1108) );
  OAI22X1TF U135 ( .A0(N634), .A1(N185), .B0(N666), .B1(N1186), .Y(N912) );
  OAI22X1TF U136 ( .A0(N680), .A1(N184), .B0(N648), .B1(N181), .Y(N1135) );
  OAI22X1TF U137 ( .A0(N163), .A1(N612), .B0(N678), .B1(N177), .Y(N1126) );
  OAI22X1TF U138 ( .A0(N618), .A1(N159), .B0(N650), .B1(N1189), .Y(N911) );
  OAI22X1TF U139 ( .A0(N694), .A1(N183), .B0(N662), .B1(N180), .Y(N1125) );
  OAI22X1TF U140 ( .A0(N690), .A1(N183), .B0(N658), .B1(N180), .Y(N1039) );
  AND2X2TF U141 ( .A(N1022), .B(N1032), .Y(N1023) );
  CLKBUFX2TF U142 ( .A(N591), .Y(N164) );
  AND2X2TF U143 ( .A(\OPER1_R1[2] ), .B(N162), .Y(N1730) );
  AND2X2TF U144 ( .A(N1033), .B(N161), .Y(N179) );
  AND2X2TF U145 ( .A(N1022), .B(N161), .Y(N182) );
  AND2X2TF U146 ( .A(N1028), .B(N161), .Y(N176) );
  NAND4X2TF U147 ( .A(N235), .B(N217), .C(N213), .D(N900), .Y(N1184) );
  AND2X2TF U148 ( .A(OPER3_R3[2]), .B(N900), .Y(N1194) );
  AND2X2TF U149 ( .A(N251), .B(N285), .Y(N1183) );
  AND2X2TF U150 ( .A(N251), .B(N262), .Y(N1181) );
  AOI32X1TF U151 ( .A0(N562), .A1(N563), .A2(N425), .B0(N561), .B1(N563), .Y(
        N591) );
  CLKINVX1TF U152 ( .A(N342), .Y(N335) );
  ADDFHX2TF U153 ( .A(N190), .B(REG_A[5]), .CI(SUB_X_292_4_N12), .CO(
        SUB_X_292_4_N11), .S(N515) );
  OAI21XLTF U154 ( .A0(N743), .A1(N742), .B0(N1198), .Y(NEXT_STATE[2]) );
  NAND3BXLTF U155 ( .AN(N897), .B(N1015), .C(N1016), .Y(N295) );
  NOR2X4TF U156 ( .A(N1016), .B(N895), .Y(N422) );
  NAND2X1TF U157 ( .A(CODE_TYPE[2]), .B(N562), .Y(N895) );
  OR2X1TF U158 ( .A(N40), .B(N781), .Y(N238) );
  CLKINVX2TF U159 ( .A(N421), .Y(N167) );
  OR2X2TF U160 ( .A(\STATE[3] ), .B(N744), .Y(N1198) );
  AND2X2TF U161 ( .A(N187), .B(N38), .Y(N838) );
  OR2X2TF U162 ( .A(N187), .B(REG_B[0]), .Y(N804) );
  NAND4XLTF U163 ( .A(N557), .B(N674), .C(N673), .D(N672), .Y(N732) );
  INVX2TF U164 ( .A(N134), .Y(N135) );
  INVX2TF U165 ( .A(N883), .Y(N136) );
  INVX2TF U166 ( .A(N838), .Y(N137) );
  INVX2TF U167 ( .A(N838), .Y(N138) );
  INVX2TF U168 ( .A(N1183), .Y(N139) );
  INVX2TF U169 ( .A(N1183), .Y(N140) );
  INVX2TF U170 ( .A(N1181), .Y(N141) );
  INVX2TF U171 ( .A(N1181), .Y(N142) );
  INVX2TF U172 ( .A(N804), .Y(N143) );
  INVX2TF U173 ( .A(N804), .Y(N144) );
  INVX2TF U174 ( .A(N1059), .Y(N145) );
  INVX2TF U175 ( .A(N1059), .Y(N146) );
  INVX2TF U176 ( .A(N1173), .Y(N147) );
  INVX2TF U177 ( .A(N1173), .Y(N148) );
  INVX2TF U178 ( .A(N858), .Y(N149) );
  INVX2TF U179 ( .A(N858), .Y(N150) );
  INVX2TF U180 ( .A(N1174), .Y(N152) );
  INVX2TF U181 ( .A(N1174), .Y(N153) );
  INVX2TF U182 ( .A(N1175), .Y(N154) );
  INVX2TF U183 ( .A(N1175), .Y(N155) );
  INVX2TF U184 ( .A(N156), .Y(N157) );
  INVX2TF U185 ( .A(N156), .Y(N158) );
  INVX2TF U186 ( .A(N1194), .Y(N159) );
  INVX2TF U187 ( .A(N1194), .Y(N160) );
  INVX2TF U188 ( .A(N1168), .Y(N161) );
  INVX2TF U189 ( .A(N1168), .Y(N162) );
  INVX2TF U190 ( .A(N1168), .Y(N163) );
  AOI22XLTF U191 ( .A0(N339), .A1(N863), .B0(N763), .B1(N861), .Y(N298) );
  NOR3X2TF U192 ( .A(N747), .B(N243), .C(\OPER1_R1[2] ), .Y(N1022) );
  AOI22X2TF U193 ( .A0(REG_C[11]), .A1(N590), .B0(N592), .B1(D_DATAIN[3]), .Y(
        N705) );
  AOI22X2TF U194 ( .A0(REG_C[10]), .A1(N590), .B0(N592), .B1(D_DATAIN[2]), .Y(
        N704) );
  AOI22X2TF U195 ( .A0(REG_C[12]), .A1(N590), .B0(N592), .B1(D_DATAIN[4]), .Y(
        N706) );
  AOI22X2TF U196 ( .A0(REG_C[8]), .A1(N590), .B0(N592), .B1(D_DATAIN[0]), .Y(
        N702) );
  AOI32X1TF U197 ( .A0(N232), .A1(N540), .A2(N741), .B0(N215), .B1(N540), .Y(
        N172) );
  NOR2BX2TF U198 ( .AN(CODE_TYPE[4]), .B(CODE_TYPE[3]), .Y(N425) );
  INVX2TF U199 ( .A(N1198), .Y(N165) );
  INVX2TF U200 ( .A(N1198), .Y(N166) );
  OAI22X2TF U201 ( .A0(N550), .A1(N564), .B0(N742), .B1(N741), .Y(N723) );
  NOR3X4TF U202 ( .A(N575), .B(N574), .C(N698), .Y(N701) );
  NOR3X4TF U203 ( .A(N575), .B(N574), .C(N576), .Y(N578) );
  NOR3X4TF U204 ( .A(N574), .B(N243), .C(N698), .Y(N697) );
  AOI22X2TF U205 ( .A0(D_ADDR[2]), .A1(N566), .B0(N565), .B1(D_DATAIN[1]), .Y(
        N581) );
  AOI22X2TF U206 ( .A0(D_ADDR[8]), .A1(N566), .B0(N565), .B1(D_DATAIN[7]), .Y(
        N588) );
  AOI22X2TF U207 ( .A0(D_ADDR[6]), .A1(N566), .B0(N565), .B1(D_DATAIN[5]), .Y(
        N585) );
  AOI22X2TF U208 ( .A0(D_ADDR[1]), .A1(N566), .B0(N565), .B1(D_DATAIN[0]), .Y(
        N580) );
  NOR3X4TF U209 ( .A(N232), .B(N745), .C(N559), .Y(N565) );
  OAI22XLTF U210 ( .A0(N639), .A1(N185), .B0(N671), .B1(N1186), .Y(N916) );
  OAI22XLTF U211 ( .A0(N633), .A1(N185), .B0(N665), .B1(N1186), .Y(N904) );
  OAI22XLTF U212 ( .A0(N617), .A1(N159), .B0(N649), .B1(N1189), .Y(N903) );
  OAI22XLTF U213 ( .A0(N623), .A1(N159), .B0(N655), .B1(N1189), .Y(N915) );
  INVX2TF U214 ( .A(N859), .Y(N168) );
  NOR2X1TF U215 ( .A(N1016), .B(N1042), .Y(N424) );
  CLKBUFX2TF U216 ( .A(N1179), .Y(N169) );
  CLKBUFX2TF U217 ( .A(N1171), .Y(N170) );
  NOR2BX2TF U218 ( .AN(N161), .B(N1030), .Y(N1171) );
  CLKBUFX2TF U219 ( .A(N1184), .Y(N171) );
  INVX2TF U220 ( .A(N1196), .Y(N1720) );
  OAI31X4TF U221 ( .A0(N1027), .A1(N1026), .A2(N1025), .B0(N1024), .Y(N1059)
         );
  NOR2X4TF U222 ( .A(N187), .B(N38), .Y(N758) );
  NOR3X4TF U223 ( .A(N875), .B(REG_B[3]), .C(N40), .Y(N870) );
  INVX2TF U224 ( .A(N1730), .Y(N1740) );
  INVX2TF U225 ( .A(N1730), .Y(N175) );
  INVX2TF U226 ( .A(N176), .Y(N177) );
  INVX2TF U227 ( .A(N176), .Y(N178) );
  INVX2TF U228 ( .A(N179), .Y(N180) );
  INVX2TF U229 ( .A(N179), .Y(N181) );
  OAI21X2TF U230 ( .A0(N896), .A1(N919), .B0(N1024), .Y(N1138) );
  OAI211X4TF U231 ( .A0(CODE_TYPE[3]), .A1(N889), .B0(N1024), .C0(N212), .Y(
        N898) );
  INVX2TF U232 ( .A(N182), .Y(N183) );
  INVX2TF U233 ( .A(N182), .Y(N184) );
  CLKBUFX2TF U234 ( .A(N1187), .Y(N185) );
  OAI22XLTF U235 ( .A0(N643), .A1(N1187), .B0(N675), .B1(N1186), .Y(N921) );
  NOR3X4TF U236 ( .A(N574), .B(N243), .C(N576), .Y(N573) );
  CLKBUFX2TF U237 ( .A(N1182), .Y(N186) );
  NOR2X1TF U238 ( .A(N258), .B(N1128), .Y(N1182) );
  AOI2BB2X2TF U239 ( .B0(D_DATAIN[6]), .B1(N592), .A0N(N418), .A1N(N164), .Y(
        N709) );
  AOI2BB2X2TF U240 ( .B0(D_DATAIN[5]), .B1(N592), .A0N(N423), .A1N(N164), .Y(
        N707) );
  AOI2BB2X2TF U241 ( .B0(D_DATAIN[7]), .B1(N592), .A0N(N416), .A1N(N164), .Y(
        N700) );
  AOI22X2TF U242 ( .A0(REG_C[9]), .A1(N590), .B0(N592), .B1(D_DATAIN[1]), .Y(
        N703) );
  NOR3X4TF U243 ( .A(N218), .B(N890), .C(N891), .Y(N592) );
  AOI22X2TF U244 ( .A0(D_ADDR[4]), .A1(N566), .B0(N565), .B1(D_DATAIN[3]), .Y(
        N583) );
  AOI22X2TF U245 ( .A0(D_ADDR[3]), .A1(N566), .B0(N565), .B1(D_DATAIN[2]), .Y(
        N582) );
  AOI22X2TF U246 ( .A0(D_ADDR[7]), .A1(N566), .B0(N565), .B1(D_DATAIN[6]), .Y(
        N586) );
  AOI22X2TF U247 ( .A0(D_ADDR[5]), .A1(N566), .B0(N565), .B1(D_DATAIN[4]), .Y(
        N584) );
  NOR3X4TF U248 ( .A(N232), .B(N215), .C(N745), .Y(N566) );
  ADDFHX2TF U249 ( .A(REG_A[15]), .B(REG_B[15]), .CI(ADD_X_292_3_N2), .CO(N492), .S(N491) );
  XOR2X1TF U250 ( .A(REG_A[0]), .B(REG_B[0]), .Y(N510) );
  NAND2BX1TF U251 ( .AN(REG_A[0]), .B(REG_B[0]), .Y(SUB_X_292_4_N16) );
  CMPR32X2TF U252 ( .A(N195), .B(REG_A[10]), .C(SUB_X_292_4_N7), .CO(
        SUB_X_292_4_N6), .S(N520) );
  CMPR32X2TF U253 ( .A(N194), .B(REG_A[9]), .C(SUB_X_292_4_N8), .CO(
        SUB_X_292_4_N7), .S(N519) );
  ADDFHX2TF U254 ( .A(N188), .B(REG_A[3]), .CI(SUB_X_292_4_N14), .CO(
        SUB_X_292_4_N13), .S(N513) );
  ADDFHX2TF U255 ( .A(N189), .B(REG_A[4]), .CI(SUB_X_292_4_N13), .CO(
        SUB_X_292_4_N12), .S(N514) );
  OAI2BB1X4TF U256 ( .A0N(N363), .A1N(N491), .B0(N308), .Y(N391) );
  AOI211X2TF U257 ( .A0(N525), .A1(N252), .B0(N307), .C0(N306), .Y(N308) );
  CLKXOR2X2TF U258 ( .A(N417), .B(N397), .Y(N389) );
  AOI21X4TF U259 ( .A0(N488), .A1(N253), .B0(N291), .Y(N417) );
  AO21X1TF U260 ( .A0(N351), .A1(N427), .B0(N136), .Y(N5140) );
  NOR2X2TF U261 ( .A(N214), .B(N218), .Y(N1044) );
  AO21X1TF U262 ( .A0(IO_DATAINA[9]), .A1(N186), .B0(N386), .Y(N474) );
  AOI21X1TF U263 ( .A0(N486), .A1(N253), .B0(N314), .Y(N397) );
  CLKBUFX2TF U264 ( .A(N363), .Y(N253) );
  CLKBUFX2TF U265 ( .A(N804), .Y(N255) );
  INVX2TF U266 ( .A(N132), .Y(N259) );
  NAND2X1TF U267 ( .A(N214), .B(N258), .Y(N891) );
  CLKBUFX2TF U268 ( .A(N421), .Y(N251) );
  NAND2X1TF U269 ( .A(N234), .B(N579), .Y(N576) );
  OAI211XLTF U270 ( .A0(N742), .A1(N211), .B0(I_ADDR[0]), .C0(N746), .Y(N554)
         );
  OAI2BB1X1TF U271 ( .A0N(N253), .A1N(N484), .B0(N362), .Y(N383) );
  NOR3X1TF U272 ( .A(N572), .B(N258), .C(N214), .Y(N889) );
  OAI211XLTF U273 ( .A0(\STATE[3] ), .A1(N741), .B0(N740), .C0(N739), .Y(
        NEXT_STATE[1]) );
  AOI31X1TF U274 ( .A0(N151), .A1(N426), .A2(N1014), .B0(N564), .Y(N738) );
  NAND2X1TF U275 ( .A(N5950), .B(N234), .Y(N698) );
  OAI2BB2X1TF U276 ( .B0(N564), .B1(N164), .A0N(N592), .A1N(N565), .Y(N579) );
  NAND2X1TF U277 ( .A(N211), .B(N557), .Y(N745) );
  AOI21X2TF U278 ( .A0(N490), .A1(N363), .B0(N294), .Y(N415) );
  CLKBUFX2TF U279 ( .A(N879), .Y(N252) );
  OR2X2TF U280 ( .A(N274), .B(N273), .Y(N363) );
  OAI21X1TF U281 ( .A0(N559), .A1(N745), .B0(N744), .Y(NEXT_STATE[3]) );
  NAND2X1TF U282 ( .A(N1024), .B(N1025), .Y(N1035) );
  NAND2X1TF U283 ( .A(N1024), .B(N1026), .Y(N1034) );
  NOR2X1TF U284 ( .A(N898), .B(N919), .Y(N900) );
  INVX2TF U285 ( .A(N1196), .Y(N1197) );
  NOR2X1TF U286 ( .A(N747), .B(N575), .Y(N1028) );
  AOI21X1TF U287 ( .A0(N563), .A1(N164), .B0(N564), .Y(N5950) );
  NOR2X2TF U288 ( .A(N232), .B(N744), .Y(N1024) );
  INVX2TF U289 ( .A(N1014), .Y(N890) );
  INVX2TF U290 ( .A(N251), .Y(N1180) );
  INVX2TF U291 ( .A(N877), .Y(N4870) );
  NOR2X2TF U292 ( .A(CODE_TYPE[3]), .B(CODE_TYPE[4]), .Y(N1014) );
  NAND2X1TF U293 ( .A(N214), .B(N218), .Y(N1021) );
  NOR2X2TF U294 ( .A(N151), .B(N572), .Y(N562) );
  NOR2X1TF U295 ( .A(N221), .B(N211), .Y(N743) );
  AOI22XLTF U296 ( .A0(REG_A[5]), .A1(N1059), .B0(IO_CONTROL[5]), .B1(N1173), 
        .Y(N1038) );
  NAND2X1TF U297 ( .A(OPER3_R3[1]), .B(N902), .Y(N1189) );
  NAND2X1TF U298 ( .A(OPER3_R3[0]), .B(N899), .Y(N1186) );
  NAND3X2TF U299 ( .A(OPER3_R3[0]), .B(OPER3_R3[1]), .C(N900), .Y(N1187) );
  NAND3X2TF U300 ( .A(N898), .B(N1138), .C(N1160), .Y(N1188) );
  NAND2X1TF U301 ( .A(N295), .B(N251), .Y(N1195) );
  NOR2X2TF U302 ( .A(N596), .B(N698), .Y(N614) );
  NOR2X2TF U303 ( .A(N596), .B(N576), .Y(N570) );
  INVX2TF U304 ( .A(N566), .Y(N564) );
  NAND3X1TF U305 ( .A(N558), .B(N215), .C(N221), .Y(N744) );
  NOR2X1TF U306 ( .A(N215), .B(\STATE[3] ), .Y(N731) );
  NAND2X2TF U307 ( .A(N880), .B(N867), .Y(N845) );
  NAND3X1TF U308 ( .A(N425), .B(N1044), .C(N251), .Y(N1128) );
  AOI21X2TF U309 ( .A0(N489), .A1(N363), .B0(N284), .Y(N419) );
  NAND3X2TF U310 ( .A(N258), .B(N1044), .C(N1014), .Y(N875) );
  NAND2X1TF U311 ( .A(N1014), .B(N889), .Y(N430) );
  NOR2X1TF U312 ( .A(N228), .B(N212), .Y(N1018) );
  OR3X1TF U313 ( .A(N562), .B(N214), .C(CODE_TYPE[3]), .Y(N560) );
  OAI211XLTF U314 ( .A0(N559), .A1(N211), .B0(N1196), .C0(N739), .Y(
        NEXT_STATE[0]) );
  AO22X1TF U315 ( .A0(N414), .A1(CF_BUF), .B0(N1195), .B1(CF), .Y(N5220) );
  AOI22XLTF U316 ( .A0(REG_A[6]), .A1(N1059), .B0(IO_CONTROL[6]), .B1(N1173), 
        .Y(N1049) );
  NOR2BX1TF U317 ( .AN(N404), .B(N1034), .Y(N1029) );
  NAND2X1TF U318 ( .A(N725), .B(I_ADDR[8]), .Y(N737) );
  NOR2X1TF U319 ( .A(N726), .B(N245), .Y(N725) );
  NOR2X2TF U320 ( .A(N564), .B(N551), .Y(N729) );
  OAI2BB2XLTF U321 ( .B0(N1197), .B1(N151), .A0N(N1197), .A1N(I_DATAIN[4]), 
        .Y(N527) );
  OAI2BB2XLTF U322 ( .B0(N1197), .B1(N212), .A0N(N1197), .A1N(I_DATAIN[7]), 
        .Y(N5240) );
  OAI2BB2XLTF U323 ( .B0(N1197), .B1(N572), .A0N(N1720), .A1N(I_DATAIN[3]), 
        .Y(N528) );
  OAI2BB2XLTF U324 ( .B0(N1197), .B1(N575), .A0N(N1720), .A1N(I_DATAIN[0]), 
        .Y(N531) );
  OAI2BB2XLTF U325 ( .B0(N1197), .B1(N574), .A0N(N1720), .A1N(I_DATAIN[1]), 
        .Y(N530) );
  OAI2BB2XLTF U326 ( .B0(N1197), .B1(N214), .A0N(N1720), .A1N(I_DATAIN[5]), 
        .Y(N526) );
  OAI2BB2XLTF U327 ( .B0(N1197), .B1(N234), .A0N(N1720), .A1N(I_DATAIN[2]), 
        .Y(N529) );
  OAI2BB2XLTF U328 ( .B0(N1197), .B1(N228), .A0N(N1720), .A1N(I_DATAIN[6]), 
        .Y(N5250) );
  NAND3X1TF U329 ( .A(N221), .B(N558), .C(N731), .Y(N1196) );
  INVX2TF U330 ( .A(N614), .Y(N597) );
  INVX2TF U331 ( .A(N697), .Y(N615) );
  INVX2TF U332 ( .A(N701), .Y(N699) );
  INVX2TF U333 ( .A(N578), .Y(N577) );
  INVX2TF U334 ( .A(N708), .Y(N710) );
  NAND2X2TF U335 ( .A(N579), .B(N1022), .Y(N567) );
  INVX2TF U336 ( .A(N573), .Y(N571) );
  INVX2TF U337 ( .A(N587), .Y(N589) );
  OAI221XLTF U338 ( .A0(REG_A[2]), .A1(N132), .B0(N225), .B1(N859), .C0(N150), 
        .Y(N798) );
  OAI221XLTF U339 ( .A0(REG_A[1]), .A1(N132), .B0(N208), .B1(N859), .C0(N150), 
        .Y(N789) );
  INVX2TF U340 ( .A(N424), .Y(N859) );
  NAND2X1TF U341 ( .A(N144), .B(REG_A[10]), .Y(N828) );
  NAND2X1TF U342 ( .A(N144), .B(REG_A[11]), .Y(N777) );
  NAND2X1TF U343 ( .A(N144), .B(REG_A[7]), .Y(N773) );
  NAND2X1TF U344 ( .A(N144), .B(REG_A[8]), .Y(N756) );
  NAND2BX1TF U345 ( .AN(N1016), .B(N264), .Y(N542) );
  NAND2X1TF U346 ( .A(N214), .B(N151), .Y(N1017) );
  NOR3X1TF U347 ( .A(N260), .B(N541), .C(N879), .Y(N543) );
  INVX2TF U348 ( .A(N1195), .Y(N414) );
  AOI211X1TF U349 ( .A0(N738), .A1(N737), .B0(N736), .C0(N735), .Y(N740) );
  OAI21X1TF U350 ( .A0(IO_CONTROL[4]), .A1(N732), .B0(N731), .Y(N733) );
  OAI21X1TF U351 ( .A0(N1179), .A1(N684), .B0(N1167), .Y(N509) );
  AOI211X1TF U352 ( .A0(IO_DATAOUTB[11]), .A1(N157), .B0(N1166), .C0(N1165), 
        .Y(N1167) );
  OAI21X1TF U353 ( .A0(N1179), .A1(N687), .B0(N1062), .Y(N458) );
  AOI211X1TF U354 ( .A0(IO_DATAOUTB[8]), .A1(N157), .B0(N1061), .C0(N1060), 
        .Y(N1062) );
  OAI21X1TF U355 ( .A0(N1179), .A1(N692), .B0(N1106), .Y(N4810) );
  AOI211X1TF U356 ( .A0(IO_DATAOUTB[3]), .A1(N158), .B0(N1105), .C0(N1104), 
        .Y(N1106) );
  OAI21X1TF U357 ( .A0(N1179), .A1(N686), .B0(N1086), .Y(N471) );
  AOI211X1TF U358 ( .A0(IO_DATAOUTB[9]), .A1(N158), .B0(N1085), .C0(N1084), 
        .Y(N1086) );
  OAI21X1TF U359 ( .A0(N1179), .A1(N681), .B0(N1114), .Y(N4850) );
  AOI211X1TF U360 ( .A0(N248), .A1(N158), .B0(N1113), .C0(N1112), .Y(N1114) );
  OAI21X1TF U361 ( .A0(N1179), .A1(N688), .B0(N1178), .Y(N5130) );
  AOI211X1TF U362 ( .A0(IO_DATAOUTB[7]), .A1(N158), .B0(N1177), .C0(N1176), 
        .Y(N1178) );
  OAI21X1TF U363 ( .A0(N169), .A1(N680), .B0(N1134), .Y(N494) );
  AOI211X1TF U364 ( .A0(N249), .A1(N157), .B0(N1133), .C0(N1132), .Y(N1134) );
  OAI21X1TF U365 ( .A0(N169), .A1(N683), .B0(N1156), .Y(N504) );
  AOI211X1TF U366 ( .A0(IO_DATAOUTB[12]), .A1(N157), .B0(N1155), .C0(N1154), 
        .Y(N1156) );
  OAI21X1TF U367 ( .A0(N169), .A1(N682), .B0(N1080), .Y(N467) );
  AOI211X1TF U368 ( .A0(N247), .A1(N157), .B0(N1079), .C0(N1078), .Y(N1080) );
  OAI21X1TF U369 ( .A0(N169), .A1(N693), .B0(N1072), .Y(N463) );
  AOI211X1TF U370 ( .A0(IO_DATAOUTB[2]), .A1(N157), .B0(N1071), .C0(N1070), 
        .Y(N1072) );
  OAI21X1TF U371 ( .A0(N169), .A1(N694), .B0(N1124), .Y(N4900) );
  AOI211X1TF U372 ( .A0(IO_DATAOUTB[1]), .A1(N157), .B0(N1123), .C0(N1122), 
        .Y(N1124) );
  OAI21X1TF U373 ( .A0(N169), .A1(N685), .B0(N1096), .Y(N4760) );
  AOI211X1TF U374 ( .A0(IO_DATAOUTB[10]), .A1(N157), .B0(N1095), .C0(N1094), 
        .Y(N1096) );
  OAI21X1TF U375 ( .A0(N631), .A1(N1740), .B0(N1148), .Y(N500) );
  AOI211X1TF U376 ( .A0(N1171), .A1(IO_DATAOUTB[0]), .B0(N1147), .C0(N1146), 
        .Y(N1148) );
  OAI21X1TF U377 ( .A0(N630), .A1(N1740), .B0(N1127), .Y(N4910) );
  AOI211X1TF U378 ( .A0(N1171), .A1(IO_DATAOUTB[1]), .B0(N1126), .C0(N1125), 
        .Y(N1127) );
  OAI21X1TF U379 ( .A0(N628), .A1(N1740), .B0(N1109), .Y(N4820) );
  AOI211X1TF U380 ( .A0(N1171), .A1(IO_DATAOUTB[3]), .B0(N1108), .C0(N1107), 
        .Y(N1109) );
  OAI21X1TF U381 ( .A0(N623), .A1(N1740), .B0(N1065), .Y(N459) );
  AOI211X1TF U382 ( .A0(N1171), .A1(IO_DATAOUTB[8]), .B0(N1064), .C0(N1063), 
        .Y(N1065) );
  OAI21X1TF U383 ( .A0(N627), .A1(N1740), .B0(N1058), .Y(N455) );
  AOI211X1TF U384 ( .A0(N1171), .A1(IO_DATAOUTB[4]), .B0(N1057), .C0(N1056), 
        .Y(N1058) );
  OAI21X1TF U385 ( .A0(N625), .A1(N1740), .B0(N1052), .Y(N451) );
  AOI211X1TF U386 ( .A0(N1171), .A1(IO_DATAOUTB[6]), .B0(N1051), .C0(N1050), 
        .Y(N1052) );
  OAI21X1TF U387 ( .A0(N626), .A1(N1740), .B0(N1041), .Y(N447) );
  AOI211X1TF U388 ( .A0(N1171), .A1(IO_DATAOUTB[5]), .B0(N1040), .C0(N1039), 
        .Y(N1041) );
  OAI22X1TF U389 ( .A0(N163), .A1(N608), .B0(N674), .B1(N178), .Y(N1040) );
  OAI21X1TF U390 ( .A0(N624), .A1(N1740), .B0(N750), .Y(N435) );
  AOI211X1TF U391 ( .A0(N170), .A1(IO_DATAOUTB[7]), .B0(N749), .C0(N748), .Y(
        N750) );
  OAI22X1TF U392 ( .A0(N162), .A1(N606), .B0(N672), .B1(N178), .Y(N749) );
  OAI21X1TF U393 ( .A0(N620), .A1(N175), .B0(N1172), .Y(N5100) );
  AOI211X1TF U394 ( .A0(N170), .A1(IO_DATAOUTB[11]), .B0(N1170), .C0(N1169), 
        .Y(N1172) );
  OAI22X1TF U395 ( .A0(N163), .A1(N602), .B0(N668), .B1(N178), .Y(N1170) );
  OAI21X1TF U396 ( .A0(N619), .A1(N175), .B0(N1159), .Y(N505) );
  AOI211X1TF U397 ( .A0(N170), .A1(IO_DATAOUTB[12]), .B0(N1158), .C0(N1157), 
        .Y(N1159) );
  OAI22X1TF U398 ( .A0(N162), .A1(N601), .B0(N667), .B1(N178), .Y(N1158) );
  OAI21X1TF U399 ( .A0(N616), .A1(N175), .B0(N1137), .Y(N495) );
  AOI211X1TF U400 ( .A0(N170), .A1(N249), .B0(N1136), .C0(N1135), .Y(N1137) );
  OAI22X1TF U401 ( .A0(N163), .A1(N598), .B0(N664), .B1(N178), .Y(N1136) );
  OAI21X1TF U402 ( .A0(N617), .A1(N175), .B0(N1117), .Y(N4860) );
  AOI211X1TF U403 ( .A0(N170), .A1(N248), .B0(N1116), .C0(N1115), .Y(N1117) );
  OAI22X1TF U404 ( .A0(N162), .A1(N599), .B0(N665), .B1(N178), .Y(N1116) );
  OAI21X1TF U405 ( .A0(N621), .A1(N175), .B0(N1099), .Y(N4770) );
  AOI211X1TF U406 ( .A0(N170), .A1(IO_DATAOUTB[10]), .B0(N1098), .C0(N1097), 
        .Y(N1099) );
  OAI22X1TF U407 ( .A0(N163), .A1(N603), .B0(N669), .B1(N178), .Y(N1098) );
  OAI21X1TF U408 ( .A0(N6220), .A1(N175), .B0(N1089), .Y(N472) );
  AOI211X1TF U409 ( .A0(N170), .A1(IO_DATAOUTB[9]), .B0(N1088), .C0(N1087), 
        .Y(N1089) );
  OAI22X1TF U410 ( .A0(N162), .A1(N604), .B0(N670), .B1(N178), .Y(N1088) );
  OAI21X1TF U411 ( .A0(N618), .A1(N175), .B0(N1083), .Y(N468) );
  AOI211X1TF U412 ( .A0(N170), .A1(N247), .B0(N1082), .C0(N1081), .Y(N1083) );
  OAI22X1TF U413 ( .A0(N163), .A1(N600), .B0(N666), .B1(N178), .Y(N1082) );
  OAI21X1TF U414 ( .A0(N629), .A1(N175), .B0(N1075), .Y(N464) );
  AOI211X1TF U415 ( .A0(N170), .A1(IO_DATAOUTB[2]), .B0(N1074), .C0(N1073), 
        .Y(N1075) );
  OAI22X1TF U416 ( .A0(N162), .A1(N611), .B0(N677), .B1(N178), .Y(N1074) );
  OAI21X1TF U417 ( .A0(N169), .A1(N695), .B0(N1145), .Y(N499) );
  AOI211X1TF U418 ( .A0(IO_DATAOUTB[0]), .A1(N158), .B0(N1144), .C0(N1143), 
        .Y(N1145) );
  OAI211X1TF U419 ( .A0(N1179), .A1(N690), .B0(N1038), .C0(N1037), .Y(N446) );
  AOI21X1TF U420 ( .A0(IO_DATAOUTB[5]), .A1(N158), .B0(N1036), .Y(N1037) );
  OAI211X1TF U421 ( .A0(N1179), .A1(N689), .B0(N1049), .C0(N1048), .Y(N450) );
  AOI21X1TF U422 ( .A0(IO_DATAOUTB[6]), .A1(N158), .B0(N1047), .Y(N1048) );
  OAI211X1TF U423 ( .A0(N1179), .A1(N691), .B0(N1055), .C0(N1054), .Y(N454) );
  AOI21X1TF U424 ( .A0(IO_DATAOUTB[4]), .A1(N158), .B0(N1053), .Y(N1054) );
  NOR2X1TF U425 ( .A(N574), .B(N243), .Y(N1033) );
  NOR2X1TF U426 ( .A(N1034), .B(N404), .Y(N1031) );
  AOI22X1TF U427 ( .A0(REG_A[4]), .A1(N1059), .B0(IO_CONTROL[4]), .B1(N1173), 
        .Y(N1055) );
  AOI31X4TF U428 ( .A0(N405), .A1(N403), .A2(N1029), .B0(N1023), .Y(N1179) );
  INVX2TF U429 ( .A(N1035), .Y(N1032) );
  OAI211X1TF U430 ( .A0(N228), .A1(N1021), .B0(N1020), .C0(N1019), .Y(N1025)
         );
  AOI32X1TF U431 ( .A0(N425), .A1(N264), .A2(N572), .B0(N1018), .B1(N1017), 
        .Y(N1020) );
  OAI21X1TF U432 ( .A0(N198), .A1(N49), .B0(N914), .Y(N441) );
  NOR3X1TF U433 ( .A(N913), .B(N912), .C(N911), .Y(N914) );
  OAI22X1TF U434 ( .A0(N682), .A1(N1184), .B0(N404), .B1(N1160), .Y(N913) );
  OAI21X1TF U435 ( .A0(N199), .A1(N1188), .B0(N906), .Y(N439) );
  NOR3X1TF U436 ( .A(N905), .B(N904), .C(N903), .Y(N906) );
  OAI22X1TF U437 ( .A0(N681), .A1(N1184), .B0(N405), .B1(N1160), .Y(N905) );
  OAI21X1TF U438 ( .A0(N193), .A1(N49), .B0(N918), .Y(N442) );
  NOR3X1TF U439 ( .A(N917), .B(N916), .C(N915), .Y(N918) );
  OAI22X1TF U440 ( .A0(N687), .A1(N1184), .B0(N235), .B1(N1160), .Y(N917) );
  OAI21X1TF U441 ( .A0(N631), .A1(N160), .B0(N1142), .Y(N498) );
  NOR3X1TF U442 ( .A(N1141), .B(N1140), .C(N1139), .Y(N1142) );
  OAI22X1TF U443 ( .A0(N663), .A1(N257), .B0(N38), .B1(N1188), .Y(N1139) );
  OAI22X1TF U444 ( .A0(N647), .A1(N1187), .B0(N679), .B1(N256), .Y(N1140) );
  OAI22X1TF U445 ( .A0(N695), .A1(N1184), .B0(N235), .B1(N1138), .Y(N1141) );
  OAI21X1TF U446 ( .A0(N630), .A1(N160), .B0(N1121), .Y(N4890) );
  NOR3X1TF U447 ( .A(N1120), .B(N1119), .C(N1118), .Y(N1121) );
  OAI22X1TF U448 ( .A0(N662), .A1(N257), .B0(N187), .B1(N1188), .Y(N1118) );
  OAI22X1TF U449 ( .A0(N646), .A1(N1187), .B0(N678), .B1(N256), .Y(N1119) );
  OAI22X1TF U450 ( .A0(N694), .A1(N1184), .B0(N217), .B1(N1138), .Y(N1120) );
  OAI21X1TF U451 ( .A0(N627), .A1(N160), .B0(N923), .Y(N443) );
  NOR3X1TF U452 ( .A(N922), .B(N921), .C(N920), .Y(N923) );
  OAI22X1TF U453 ( .A0(N659), .A1(N257), .B0(N189), .B1(N1188), .Y(N920) );
  OAI22X1TF U454 ( .A0(N691), .A1(N171), .B0(N403), .B1(N1185), .Y(N922) );
  OAI21X1TF U455 ( .A0(N626), .A1(N160), .B0(N1013), .Y(N445) );
  NOR3X1TF U456 ( .A(N1012), .B(N1011), .C(N1010), .Y(N1013) );
  OAI22X1TF U457 ( .A0(N658), .A1(N257), .B0(N190), .B1(N1188), .Y(N1010) );
  OAI22X1TF U458 ( .A0(N642), .A1(N1187), .B0(N674), .B1(N256), .Y(N1011) );
  OAI22X1TF U459 ( .A0(N690), .A1(N171), .B0(N404), .B1(N1185), .Y(N1012) );
  OAI21X1TF U460 ( .A0(N625), .A1(N160), .B0(N1009), .Y(N444) );
  NOR3X1TF U461 ( .A(N926), .B(N925), .C(N924), .Y(N1009) );
  OAI22X1TF U462 ( .A0(N657), .A1(N257), .B0(N191), .B1(N1188), .Y(N924) );
  OAI22X1TF U463 ( .A0(N641), .A1(N1187), .B0(N673), .B1(N256), .Y(N925) );
  OAI22X1TF U464 ( .A0(N689), .A1(N171), .B0(N405), .B1(N1185), .Y(N926) );
  OAI21X1TF U465 ( .A0(N624), .A1(N160), .B0(N1193), .Y(N5160) );
  NOR3X1TF U466 ( .A(N1192), .B(N1191), .C(N1190), .Y(N1193) );
  OAI22X1TF U467 ( .A0(N656), .A1(N257), .B0(N192), .B1(N1188), .Y(N1190) );
  OAI22X1TF U468 ( .A0(N640), .A1(N1187), .B0(N672), .B1(N256), .Y(N1191) );
  OAI22X1TF U469 ( .A0(N406), .A1(N1185), .B0(N688), .B1(N1184), .Y(N1192) );
  OAI21X1TF U470 ( .A0(N628), .A1(N160), .B0(N1103), .Y(N4800) );
  NOR3X1TF U471 ( .A(N1102), .B(N1101), .C(N1100), .Y(N1103) );
  OAI22X1TF U472 ( .A0(N660), .A1(N257), .B0(N188), .B1(N1188), .Y(N1100) );
  OAI22X1TF U473 ( .A0(N644), .A1(N1187), .B0(N676), .B1(N256), .Y(N1101) );
  OAI22X1TF U474 ( .A0(N692), .A1(N1184), .B0(N402), .B1(N1138), .Y(N1102) );
  OAI21X1TF U475 ( .A0(N196), .A1(N49), .B0(N1164), .Y(N508) );
  NOR3X1TF U476 ( .A(N1163), .B(N1162), .C(N1161), .Y(N1164) );
  OAI22X1TF U477 ( .A0(N620), .A1(N159), .B0(N652), .B1(N1189), .Y(N1161) );
  OAI22X1TF U478 ( .A0(N636), .A1(N185), .B0(N668), .B1(N256), .Y(N1162) );
  OAI22X1TF U479 ( .A0(N684), .A1(N171), .B0(N402), .B1(N1160), .Y(N1163) );
  OAI21X1TF U480 ( .A0(N197), .A1(N49), .B0(N1153), .Y(N503) );
  NOR3X1TF U481 ( .A(N1152), .B(N1151), .C(N1150), .Y(N1153) );
  OAI22X1TF U482 ( .A0(N619), .A1(N159), .B0(N651), .B1(N1189), .Y(N1150) );
  OAI22X1TF U483 ( .A0(N635), .A1(N185), .B0(N667), .B1(N256), .Y(N1151) );
  OAI22X1TF U484 ( .A0(N683), .A1(N171), .B0(N403), .B1(N1160), .Y(N1152) );
  OAI21X1TF U485 ( .A0(N629), .A1(N160), .B0(N1069), .Y(N462) );
  NOR3X1TF U486 ( .A(N1068), .B(N1067), .C(N1066), .Y(N1069) );
  OAI22X1TF U487 ( .A0(N661), .A1(N257), .B0(N133), .B1(N1188), .Y(N1066) );
  OAI22X1TF U488 ( .A0(N645), .A1(N185), .B0(N677), .B1(N256), .Y(N1067) );
  OAI22X1TF U489 ( .A0(N693), .A1(N1184), .B0(N213), .B1(N1138), .Y(N1068) );
  OAI21X1TF U490 ( .A0(N194), .A1(N49), .B0(N910), .Y(N440) );
  NOR3X1TF U491 ( .A(N909), .B(N908), .C(N907), .Y(N910) );
  OAI22X1TF U492 ( .A0(N6220), .A1(N159), .B0(N654), .B1(N257), .Y(N907) );
  OAI22X1TF U493 ( .A0(N686), .A1(N171), .B0(N217), .B1(N1160), .Y(N909) );
  OAI21X1TF U494 ( .A0(N195), .A1(N49), .B0(N1093), .Y(N475) );
  NOR3X1TF U495 ( .A(N1092), .B(N1091), .C(N1090), .Y(N1093) );
  OAI22X1TF U496 ( .A0(N621), .A1(N159), .B0(N653), .B1(N257), .Y(N1090) );
  NOR2X1TF U497 ( .A(OPER3_R3[0]), .B(N901), .Y(N902) );
  OAI22X1TF U498 ( .A0(N637), .A1(N1187), .B0(N669), .B1(N256), .Y(N1091) );
  NOR2X1TF U499 ( .A(OPER3_R3[1]), .B(N901), .Y(N899) );
  OAI22X1TF U500 ( .A0(N685), .A1(N171), .B0(N213), .B1(N1160), .Y(N1092) );
  NAND2X2TF U501 ( .A(N897), .B(N1024), .Y(N1160) );
  OAI211X1TF U502 ( .A0(N895), .A1(N212), .B0(N894), .C0(N893), .Y(N919) );
  INVX2TF U503 ( .A(N1021), .Y(N426) );
  AOI21X1TF U504 ( .A0(N892), .A1(N891), .B0(N890), .Y(N896) );
  AOI211X1TF U505 ( .A0(N752), .A1(N751), .B0(CODE_TYPE[2]), .C0(N1043), .Y(
        N897) );
  AOI21X1TF U506 ( .A0(D_ADDR[2]), .A1(N729), .B0(N712), .Y(N816) );
  OAI21X1TF U507 ( .A0(N723), .A1(N241), .B0(N711), .Y(N712) );
  OAI211X1TF U508 ( .A0(I_ADDR[1]), .A1(I_ADDR[2]), .B0(N720), .C0(N713), .Y(
        N711) );
  AOI211X1TF U509 ( .A0(N729), .A1(D_ADDR[3]), .B0(N715), .C0(N714), .Y(N815)
         );
  AOI211X1TF U510 ( .A0(N713), .A1(N216), .B0(N716), .C0(N724), .Y(N714) );
  NOR2X1TF U511 ( .A(N216), .B(N723), .Y(N715) );
  AOI21X1TF U512 ( .A0(D_ADDR[1]), .A1(N729), .B0(N552), .Y(N865) );
  AOI22X1TF U513 ( .A0(I_ADDR[1]), .A1(N723), .B0(N724), .B1(N233), .Y(N552)
         );
  AOI211X1TF U514 ( .A0(N729), .A1(D_ADDR[7]), .B0(N728), .C0(N727), .Y(N808)
         );
  AOI211X1TF U515 ( .A0(N726), .A1(N245), .B0(N725), .C0(N724), .Y(N727) );
  NOR2X1TF U516 ( .A(N245), .B(N723), .Y(N728) );
  AOI211X1TF U517 ( .A0(N729), .A1(D_ADDR[5]), .B0(N719), .C0(N718), .Y(N813)
         );
  AOI211X1TF U518 ( .A0(N717), .A1(N242), .B0(N721), .C0(N724), .Y(N718) );
  NOR2X1TF U519 ( .A(N242), .B(N723), .Y(N719) );
  OAI32X1TF U520 ( .A0(N553), .A1(N725), .A2(I_ADDR[8]), .B0(N720), .B1(N553), 
        .Y(N864) );
  INVX2TF U521 ( .A(N724), .Y(N720) );
  INVX2TF U522 ( .A(N723), .Y(N722) );
  NOR2X1TF U523 ( .A(N717), .B(N242), .Y(N721) );
  NOR3X1TF U524 ( .A(N233), .B(N241), .C(N216), .Y(N716) );
  AOI32X1TF U525 ( .A0(N549), .A1(N1018), .A2(N244), .B0(N548), .B1(N1018), 
        .Y(N551) );
  OAI22X1TF U526 ( .A0(N751), .A1(N244), .B0(N547), .B1(N546), .Y(N548) );
  OAI22X1TF U527 ( .A0(CF), .A1(N892), .B0(N545), .B1(N214), .Y(N546) );
  AOI21X1TF U528 ( .A0(CF), .A1(N218), .B0(N151), .Y(N545) );
  AOI22X1TF U529 ( .A0(N697), .A1(N707), .B0(N650), .B1(N615), .Y(N944) );
  AOI22X1TF U530 ( .A0(N614), .A1(N707), .B0(N666), .B1(N597), .Y(N952) );
  AOI22X1TF U531 ( .A0(N701), .A1(N707), .B0(N634), .B1(N699), .Y(N936) );
  AOI22X1TF U532 ( .A0(N697), .A1(N700), .B0(N648), .B1(N615), .Y(N942) );
  AOI22X1TF U533 ( .A0(N701), .A1(N700), .B0(N632), .B1(N699), .Y(N934) );
  AOI22X1TF U534 ( .A0(N614), .A1(N700), .B0(N664), .B1(N597), .Y(N950) );
  AOI22X1TF U535 ( .A0(N701), .A1(N709), .B0(N633), .B1(N699), .Y(N935) );
  AOI22X1TF U536 ( .A0(N697), .A1(N709), .B0(N649), .B1(N615), .Y(N943) );
  AOI22X1TF U537 ( .A0(N614), .A1(N709), .B0(N665), .B1(N597), .Y(N951) );
  AOI22X1TF U538 ( .A0(N710), .A1(N700), .B0(N616), .B1(N708), .Y(N1006) );
  AOI22X1TF U539 ( .A0(N710), .A1(N707), .B0(N618), .B1(N708), .Y(N928) );
  AOI22X1TF U540 ( .A0(N710), .A1(N709), .B0(N617), .B1(N708), .Y(N927) );
  AOI22X1TF U541 ( .A0(N5940), .A1(N709), .B0(N681), .B1(N593), .Y(N959) );
  AOI22X1TF U542 ( .A0(N5940), .A1(N707), .B0(N682), .B1(N593), .Y(N960) );
  AOI22X1TF U543 ( .A0(N5940), .A1(N700), .B0(N680), .B1(N593), .Y(N958) );
  AOI22X1TF U544 ( .A0(N578), .A1(N583), .B0(N644), .B1(N577), .Y(N978) );
  AOI22X1TF U545 ( .A0(N578), .A1(N588), .B0(N640), .B1(N577), .Y(N974) );
  AOI22X1TF U546 ( .A0(N570), .A1(N583), .B0(N676), .B1(N569), .Y(N994) );
  AOI22X1TF U547 ( .A0(N570), .A1(N582), .B0(N677), .B1(N569), .Y(N995) );
  AOI22X1TF U548 ( .A0(N614), .A1(N703), .B0(N670), .B1(N597), .Y(N956) );
  AOI22X1TF U549 ( .A0(N614), .A1(N705), .B0(N668), .B1(N597), .Y(N954) );
  AOI22X1TF U550 ( .A0(N570), .A1(N584), .B0(N675), .B1(N569), .Y(N993) );
  AOI22X1TF U552 ( .A0(N578), .A1(N586), .B0(N641), .B1(N577), .Y(N975) );
  AOI22X1TF U553 ( .A0(N578), .A1(N582), .B0(N645), .B1(N577), .Y(N979) );
  AOI22X1TF U554 ( .A0(N570), .A1(N588), .B0(N672), .B1(N569), .Y(N990) );
  AOI22X1TF U555 ( .A0(N570), .A1(N586), .B0(N673), .B1(N569), .Y(N991) );
  AOI22X1TF U556 ( .A0(N570), .A1(N585), .B0(N674), .B1(N569), .Y(N992) );
  AOI22X1TF U557 ( .A0(N697), .A1(N703), .B0(N654), .B1(N615), .Y(N948) );
  AOI22X1TF U558 ( .A0(N578), .A1(N581), .B0(N646), .B1(N577), .Y(N980) );
  AOI22X1TF U559 ( .A0(N570), .A1(N580), .B0(N679), .B1(N569), .Y(N997) );
  AOI22X1TF U560 ( .A0(N701), .A1(N703), .B0(N638), .B1(N699), .Y(N940) );
  AOI22X1TF U561 ( .A0(N578), .A1(N584), .B0(N643), .B1(N577), .Y(N977) );
  AOI22X1TF U562 ( .A0(N578), .A1(N580), .B0(N647), .B1(N577), .Y(N981) );
  AOI22X1TF U563 ( .A0(N578), .A1(N585), .B0(N642), .B1(N577), .Y(N976) );
  AOI22X1TF U564 ( .A0(N570), .A1(N581), .B0(N678), .B1(N569), .Y(N996) );
  INVX2TF U565 ( .A(N570), .Y(N569) );
  AOI22X1TF U566 ( .A0(N710), .A1(N706), .B0(N619), .B1(N708), .Y(N929) );
  AOI22X1TF U567 ( .A0(N710), .A1(N702), .B0(N623), .B1(N708), .Y(N933) );
  AOI22X1TF U568 ( .A0(N710), .A1(N703), .B0(N6220), .B1(N708), .Y(N932) );
  AOI22X1TF U569 ( .A0(N710), .A1(N705), .B0(N620), .B1(N708), .Y(N930) );
  AOI22X1TF U570 ( .A0(N710), .A1(N704), .B0(N621), .B1(N708), .Y(N931) );
  NAND4X2TF U571 ( .A(N575), .B(N574), .C(\OPER1_R1[2] ), .D(N5950), .Y(N708)
         );
  AOI22X1TF U572 ( .A0(N5940), .A1(N703), .B0(N686), .B1(N593), .Y(N964) );
  AOI22X1TF U573 ( .A0(N5940), .A1(N705), .B0(N684), .B1(N593), .Y(N962) );
  AOI22X1TF U574 ( .A0(N5940), .A1(N704), .B0(N685), .B1(N593), .Y(N963) );
  AOI22X1TF U575 ( .A0(N5940), .A1(N706), .B0(N683), .B1(N593), .Y(N961) );
  AOI22X1TF U576 ( .A0(N5940), .A1(N702), .B0(N687), .B1(N593), .Y(N965) );
  INVX2TF U577 ( .A(N164), .Y(N590) );
  NAND2X2TF U578 ( .A(N5950), .B(N1022), .Y(N593) );
  AOI22X1TF U579 ( .A0(N568), .A1(N584), .B0(N691), .B1(N567), .Y(N1001) );
  AOI22X1TF U580 ( .A0(N568), .A1(N585), .B0(N690), .B1(N567), .Y(N1000) );
  AOI22X1TF U581 ( .A0(N568), .A1(N582), .B0(N693), .B1(N567), .Y(N1003) );
  AOI22X1TF U582 ( .A0(N568), .A1(N583), .B0(N692), .B1(N567), .Y(N1002) );
  AOI22X1TF U583 ( .A0(N568), .A1(N586), .B0(N689), .B1(N567), .Y(N999) );
  AOI22X1TF U584 ( .A0(N568), .A1(N580), .B0(N695), .B1(N567), .Y(N1005) );
  AOI22X1TF U585 ( .A0(N568), .A1(N581), .B0(N694), .B1(N567), .Y(N1004) );
  AOI22X1TF U586 ( .A0(N568), .A1(N588), .B0(N688), .B1(N567), .Y(N998) );
  INVX2TF U587 ( .A(N567), .Y(N568) );
  AOI22X1TF U588 ( .A0(N573), .A1(N583), .B0(N660), .B1(N571), .Y(N986) );
  AOI22X1TF U589 ( .A0(N573), .A1(N584), .B0(N659), .B1(N571), .Y(N985) );
  AOI22X1TF U590 ( .A0(N573), .A1(N582), .B0(N661), .B1(N571), .Y(N987) );
  AOI22X1TF U591 ( .A0(N573), .A1(N580), .B0(N663), .B1(N571), .Y(N989) );
  AOI22X1TF U592 ( .A0(N573), .A1(N586), .B0(N657), .B1(N571), .Y(N983) );
  AOI22X1TF U593 ( .A0(N589), .A1(N583), .B0(N628), .B1(N587), .Y(N970) );
  AOI22X1TF U594 ( .A0(N589), .A1(N582), .B0(N629), .B1(N587), .Y(N971) );
  AOI22X1TF U595 ( .A0(N589), .A1(N586), .B0(N625), .B1(N587), .Y(N967) );
  AOI22X1TF U596 ( .A0(N589), .A1(N584), .B0(N627), .B1(N587), .Y(N969) );
  AOI22X1TF U597 ( .A0(N589), .A1(N580), .B0(N631), .B1(N587), .Y(N973) );
  AOI22X1TF U598 ( .A0(N589), .A1(N581), .B0(N630), .B1(N587), .Y(N972) );
  AOI22X1TF U599 ( .A0(N589), .A1(N588), .B0(N624), .B1(N587), .Y(N966) );
  AOI22X1TF U600 ( .A0(N589), .A1(N585), .B0(N626), .B1(N587), .Y(N968) );
  NAND4X2TF U601 ( .A(N574), .B(N575), .C(\OPER1_R1[2] ), .D(N579), .Y(N587)
         );
  INVX2TF U602 ( .A(N592), .Y(N563) );
  OAI32X1TF U603 ( .A0(N696), .A1(N1024), .A2(N250), .B0(N555), .B1(N696), .Y(
        N1007) );
  AOI22X1TF U604 ( .A0(I_ADDR[0]), .A1(N598), .B0(N606), .B1(N230), .Y(
        D_DATAOUT[7]) );
  AOI22X1TF U605 ( .A0(I_ADDR[0]), .A1(N599), .B0(N607), .B1(N230), .Y(
        D_DATAOUT[6]) );
  AOI22X1TF U606 ( .A0(I_ADDR[0]), .A1(N600), .B0(N608), .B1(N230), .Y(
        D_DATAOUT[5]) );
  AOI22X1TF U607 ( .A0(I_ADDR[0]), .A1(N601), .B0(N609), .B1(N230), .Y(
        D_DATAOUT[4]) );
  AOI22X1TF U608 ( .A0(I_ADDR[0]), .A1(N602), .B0(N610), .B1(N230), .Y(
        D_DATAOUT[3]) );
  AOI22X1TF U609 ( .A0(I_ADDR[0]), .A1(N603), .B0(N611), .B1(N230), .Y(
        D_DATAOUT[2]) );
  AOI22X1TF U610 ( .A0(I_ADDR[0]), .A1(N604), .B0(N612), .B1(N230), .Y(
        D_DATAOUT[1]) );
  AOI22X1TF U611 ( .A0(I_ADDR[0]), .A1(N605), .B0(N613), .B1(N230), .Y(
        D_DATAOUT[0]) );
  OAI211X1TF U612 ( .A0(N730), .A1(N554), .B0(N734), .C0(N555), .Y(N1008) );
  NOR2X1TF U613 ( .A(N251), .B(N565), .Y(N734) );
  INVX2TF U614 ( .A(N1024), .Y(N746) );
  INVX2TF U615 ( .A(N731), .Y(N742) );
  INVX2TF U616 ( .A(N745), .Y(N730) );
  AOI21X1TF U617 ( .A0(N378), .A1(N1183), .B0(N377), .Y(N379) );
  AOI22X1TF U618 ( .A0(N254), .A1(IO_DATAINB[4]), .B0(D_ADDR[5]), .B1(N1180), 
        .Y(N375) );
  AOI22X1TF U619 ( .A0(N1149), .A1(IO_STATUS[1]), .B0(N186), .B1(IO_DATAINA[1]), .Y(N1130) );
  AOI22X1TF U620 ( .A0(IO_DATAINB[1]), .A1(N409), .B0(D_ADDR[2]), .B1(N167), 
        .Y(N1131) );
  AOI21X1TF U621 ( .A0(N383), .A1(N1181), .B0(N381), .Y(N382) );
  OAI21X1TF U622 ( .A0(N400), .A1(N139), .B0(N380), .Y(N381) );
  AOI22X1TF U623 ( .A0(N254), .A1(IO_DATAINB[8]), .B0(REG_C[8]), .B1(N1180), 
        .Y(N380) );
  OAI211X1TF U624 ( .A0(N387), .A1(N141), .B0(N385), .C0(N384), .Y(N386) );
  AOI21X1TF U625 ( .A0(N518), .A1(N252), .B0(N361), .Y(N362) );
  OAI21X1TF U626 ( .A0(N843), .A1(N833), .B0(N360), .Y(N361) );
  OAI22X1TF U627 ( .A0(N846), .A1(N848), .B0(N836), .B1(N885), .Y(N358) );
  OAI22X1TF U628 ( .A0(N837), .A1(N845), .B0(N844), .B1(N878), .Y(N835) );
  NOR2X1TF U629 ( .A(N357), .B(N239), .Y(N359) );
  AOI22X1TF U630 ( .A0(REG_A[8]), .A1(N424), .B0(N422), .B1(N239), .Y(N831) );
  AOI22X1TF U631 ( .A0(N254), .A1(IO_DATAINB[9]), .B0(REG_C[9]), .B1(N1180), 
        .Y(N385) );
  AOI21X1TF U632 ( .A0(N485), .A1(N253), .B0(N320), .Y(N387) );
  AOI211X1TF U633 ( .A0(REG_A[9]), .A1(N318), .B0(N825), .C0(N317), .Y(N319)
         );
  OAI21X1TF U634 ( .A0(N823), .A1(N843), .B0(N316), .Y(N317) );
  AOI211X1TF U635 ( .A0(N870), .A1(N853), .B0(N315), .C0(N826), .Y(N316) );
  OAI22X1TF U636 ( .A0(N852), .A1(N845), .B0(N821), .B1(N238), .Y(N826) );
  NOR2X1TF U637 ( .A(N878), .B(N824), .Y(N315) );
  AOI22X1TF U638 ( .A0(REG_A[9]), .A1(N168), .B0(N260), .B1(N220), .Y(N822) );
  OAI211X1TF U639 ( .A0(N410), .A1(N142), .B0(N1046), .C0(N1045), .Y(N449) );
  AOI22X1TF U640 ( .A0(IO_DATAINA[5]), .A1(N186), .B0(N1183), .B1(N376), .Y(
        N1045) );
  OR2X2TF U641 ( .A(N847), .B(N356), .Y(N376) );
  AOI22X1TF U642 ( .A0(N480), .A1(N363), .B0(N879), .B1(N514), .Y(N349) );
  OAI22X1TF U643 ( .A0(N837), .A1(N851), .B0(N878), .B1(N836), .Y(N849) );
  INVX2TF U644 ( .A(N832), .Y(N836) );
  INVX2TF U645 ( .A(N862), .Y(N837) );
  INVX2TF U646 ( .A(N866), .Y(N846) );
  AOI22X1TF U647 ( .A0(REG_A[4]), .A1(N168), .B0(N422), .B1(N237), .Y(N842) );
  AOI22X1TF U648 ( .A0(IO_DATAINB[5]), .A1(N409), .B0(D_ADDR[6]), .B1(N167), 
        .Y(N1046) );
  AOI21X1TF U649 ( .A0(N407), .A1(N1183), .B0(N401), .Y(N408) );
  OAI21X1TF U650 ( .A0(N400), .A1(N141), .B0(N399), .Y(N401) );
  AOI22X1TF U651 ( .A0(N409), .A1(IO_DATAINB[7]), .B0(D_ADDR[8]), .B1(N1180), 
        .Y(N399) );
  OAI211X1TF U652 ( .A0(N411), .A1(N140), .B0(N1111), .C0(N1110), .Y(N4840) );
  AOI22X1TF U653 ( .A0(IO_DATAINA[3]), .A1(N186), .B0(N1181), .B1(N378), .Y(
        N1110) );
  OAI211X1TF U654 ( .A0(N820), .A1(N851), .B0(N819), .C0(N367), .Y(N378) );
  OAI21X1TF U655 ( .A0(N806), .A1(N843), .B0(N365), .Y(N366) );
  AOI21X1TF U656 ( .A0(N513), .A1(N879), .B0(N364), .Y(N365) );
  AOI211X1TF U657 ( .A0(REG_A[5]), .A1(N144), .B0(N803), .C0(N802), .Y(N805)
         );
  INVX2TF U658 ( .A(N763), .Y(N806) );
  NOR4BX1TF U659 ( .AN(N767), .B(N766), .C(N765), .D(N764), .Y(N807) );
  AOI221X1TF U660 ( .A0(N219), .A1(N422), .B0(REG_A[3]), .B1(N168), .C0(N811), 
        .Y(N817) );
  OAI21X1TF U661 ( .A0(REG_B[3]), .A1(N132), .B0(N809), .Y(N818) );
  AOI211X1TF U662 ( .A0(REG_A[11]), .A1(N427), .B0(N770), .C0(N769), .Y(N820)
         );
  OAI22X1TF U663 ( .A0(N785), .A1(N210), .B0(N255), .B1(N226), .Y(N769) );
  INVX2TF U664 ( .A(N768), .Y(N770) );
  AOI22X1TF U665 ( .A0(IO_DATAINB[3]), .A1(N409), .B0(D_ADDR[4]), .B1(N1180), 
        .Y(N1111) );
  AOI21X1TF U666 ( .A0(N407), .A1(N1181), .B0(N373), .Y(N374) );
  OAI21X1TF U667 ( .A0(N410), .A1(N140), .B0(N372), .Y(N373) );
  AOI22X1TF U668 ( .A0(N254), .A1(IO_DATAINB[6]), .B0(D_ADDR[7]), .B1(N1180), 
        .Y(N372) );
  AOI211X1TF U669 ( .A0(N481), .A1(N253), .B0(N338), .C0(N337), .Y(N410) );
  AOI211X1TF U670 ( .A0(N855), .A1(N335), .B0(N856), .C0(N334), .Y(N336) );
  OAI22X1TF U671 ( .A0(N852), .A1(N851), .B0(N850), .B1(N209), .Y(N856) );
  OAI21X1TF U672 ( .A0(N843), .A1(N877), .B0(N326), .Y(N407) );
  AOI211X1TF U673 ( .A0(N482), .A1(N363), .B0(N325), .C0(N761), .Y(N326) );
  AOI22X1TF U674 ( .A0(REG_A[6]), .A1(N168), .B0(N260), .B1(N240), .Y(N757) );
  OAI211X1TF U675 ( .A0(N324), .A1(N240), .B0(N323), .C0(N322), .Y(N325) );
  AOI211X1TF U676 ( .A0(N854), .A1(N793), .B0(N321), .C0(N762), .Y(N322) );
  OAI22X1TF U677 ( .A0(N886), .A1(N878), .B0(N753), .B1(N795), .Y(N762) );
  NOR2X1TF U678 ( .A(N848), .B(N790), .Y(N321) );
  OAI211X1TF U679 ( .A0(N413), .A1(N140), .B0(N1077), .C0(N1076), .Y(N466) );
  INVX2TF U680 ( .A(N370), .Y(N411) );
  OAI211X1TF U681 ( .A0(N886), .A1(N843), .B0(N799), .C0(N341), .Y(N370) );
  AOI211X1TF U682 ( .A0(N512), .A1(N879), .B0(N800), .C0(N340), .Y(N341) );
  INVX2TF U683 ( .A(N845), .Y(N854) );
  INVX2TF U684 ( .A(N790), .Y(N801) );
  OAI22X1TF U685 ( .A0(N796), .A1(N848), .B0(N881), .B1(N795), .Y(N800) );
  AOI211X1TF U686 ( .A0(REG_A[4]), .A1(N144), .B0(N792), .C0(N791), .Y(N796)
         );
  AOI22X1TF U687 ( .A0(N135), .A1(N798), .B0(REG_A[2]), .B1(N797), .Y(N799) );
  OAI21X1TF U688 ( .A0(N135), .A1(N132), .B0(N809), .Y(N797) );
  AOI22X1TF U689 ( .A0(IO_DATAINB[2]), .A1(N409), .B0(D_ADDR[3]), .B1(N167), 
        .Y(N1077) );
  INVX2TF U690 ( .A(N371), .Y(N413) );
  AOI21X1TF U691 ( .A0(N477), .A1(N253), .B0(N343), .Y(N345) );
  OAI211X1TF U692 ( .A0(N237), .A1(N785), .B0(N784), .C0(N783), .Y(N786) );
  OAI32X1TF U693 ( .A0(N208), .A1(REG_B[1]), .A2(N132), .B0(N809), .B1(N208), 
        .Y(N788) );
  INVX2TF U694 ( .A(N852), .Y(N780) );
  AOI21X1TF U695 ( .A0(IO_DATAINA[0]), .A1(N186), .B0(N394), .Y(N395) );
  OAI211X1TF U696 ( .A0(N412), .A1(N141), .B0(N393), .C0(N392), .Y(N394) );
  NOR2X1TF U697 ( .A(N39), .B(N1128), .Y(N1149) );
  AOI22X1TF U698 ( .A0(N254), .A1(IO_DATAINB[0]), .B0(D_ADDR[1]), .B1(N1180), 
        .Y(N393) );
  AND2X2TF U699 ( .A(N251), .B(N369), .Y(N409) );
  AND2X2TF U700 ( .A(N425), .B(N368), .Y(N369) );
  INVX2TF U701 ( .A(N1042), .Y(N368) );
  AOI211X1TF U702 ( .A0(REG_A[0]), .A1(N332), .B0(N331), .C0(N330), .Y(N412)
         );
  OAI211X1TF U703 ( .A0(N875), .A1(N876), .B0(N874), .C0(N329), .Y(N330) );
  AOI22X1TF U704 ( .A0(N252), .A1(N510), .B0(N476), .B1(N253), .Y(N329) );
  OAI31X1TF U705 ( .A0(N873), .A1(N872), .A2(N871), .B0(N870), .Y(N874) );
  NOR2X1TF U706 ( .A(N255), .B(N225), .Y(N871) );
  NOR2X1TF U707 ( .A(N869), .B(N208), .Y(N872) );
  OAI22X1TF U708 ( .A0(REG_A[0]), .A1(N132), .B0(N859), .B1(N222), .Y(N328) );
  OAI21X1TF U709 ( .A0(REG_B[0]), .A1(N132), .B0(N327), .Y(N332) );
  OAI211X1TF U710 ( .A0(N877), .A1(N878), .B0(N313), .C0(N312), .Y(N314) );
  NOR3X1TF U711 ( .A(N311), .B(N887), .C(N310), .Y(N312) );
  AOI22X1TF U712 ( .A0(N40), .A1(N794), .B0(N793), .B1(N133), .Y(N881) );
  OAI211X1TF U713 ( .A0(N138), .A1(N223), .B0(N760), .C0(N759), .Y(N793) );
  INVX2TF U714 ( .A(N875), .Y(N880) );
  OAI22X1TF U715 ( .A0(N886), .A1(N885), .B0(N884), .B1(N223), .Y(N887) );
  OAI211X1TF U716 ( .A0(N452), .A1(N197), .B0(N290), .C0(N289), .Y(N291) );
  AOI211X1TF U717 ( .A0(REG_A[12]), .A1(N288), .B0(N287), .C0(N286), .Y(N289)
         );
  OAI211X1TF U718 ( .A0(N227), .A1(N138), .B0(N460), .C0(N432), .Y(N862) );
  OAI211X1TF U719 ( .A0(N220), .A1(N785), .B0(N760), .C0(N828), .Y(N431) );
  NOR2X1TF U720 ( .A(N782), .B(N456), .Y(N287) );
  INVX2TF U721 ( .A(N844), .Y(N434) );
  AOI211X1TF U722 ( .A0(REG_A[4]), .A1(N427), .B0(N792), .C0(N433), .Y(N844)
         );
  OAI22X1TF U723 ( .A0(N785), .A1(N208), .B0(N255), .B1(N225), .Y(N433) );
  NOR2X1TF U724 ( .A(N869), .B(N219), .Y(N792) );
  NOR2X1TF U725 ( .A(N138), .B(N222), .Y(N832) );
  INVX2TF U726 ( .A(N833), .Y(N448) );
  NOR4X1TF U727 ( .A(N754), .B(N791), .C(N830), .D(N839), .Y(N833) );
  NOR2X1TF U728 ( .A(N240), .B(N255), .Y(N839) );
  NOR2X1TF U729 ( .A(N137), .B(N239), .Y(N830) );
  NOR2X1TF U730 ( .A(N785), .B(N209), .Y(N791) );
  NOR2X1TF U731 ( .A(N869), .B(N224), .Y(N754) );
  INVX2TF U732 ( .A(N132), .Y(N260) );
  AOI211X1TF U733 ( .A0(REG_A[13]), .A1(N282), .B0(N281), .C0(N280), .Y(N283)
         );
  OAI21X1TF U734 ( .A0(N852), .A1(N848), .B0(N279), .Y(N280) );
  AOI211X1TF U735 ( .A0(N278), .A1(N855), .B0(N277), .C0(N276), .Y(N279) );
  AOI31X1TF U736 ( .A0(N777), .A1(N768), .A2(N767), .B0(N843), .Y(N276) );
  NOR2X1TF U737 ( .A(N878), .B(N823), .Y(N277) );
  NOR4BBX1TF U738 ( .AN(N773), .BN(N778), .C(N764), .D(N802), .Y(N823) );
  NOR2X1TF U739 ( .A(N240), .B(N785), .Y(N802) );
  NOR2X1TF U740 ( .A(N239), .B(N869), .Y(N764) );
  OAI22X1TF U741 ( .A0(N133), .A1(N781), .B0(N824), .B1(N40), .Y(N855) );
  AOI211X1TF U742 ( .A0(REG_A[2]), .A1(N758), .B0(N428), .C0(N803), .Y(N824)
         );
  NOR2X1TF U743 ( .A(N869), .B(N237), .Y(N803) );
  OAI22X1TF U744 ( .A0(N138), .A1(N209), .B0(N255), .B1(N219), .Y(N428) );
  INVX2TF U745 ( .A(N821), .Y(N278) );
  AOI21X1TF U746 ( .A0(N427), .A1(REG_A[13]), .B0(N429), .Y(N852) );
  OAI22X1TF U747 ( .A0(N255), .A1(N229), .B0(N869), .B1(N210), .Y(N429) );
  NOR4BX1TF U748 ( .AN(N5110), .B(N501), .C(N506), .D(N292), .Y(N293) );
  NOR3X1TF U749 ( .A(N753), .B(REG_B[3]), .C(N875), .Y(N292) );
  AOI221X1TF U750 ( .A0(REG_B[0]), .A1(N229), .B0(N38), .B1(N210), .C0(
        REG_B[1]), .Y(N794) );
  AOI31X1TF U751 ( .A0(N465), .A1(N827), .A2(N460), .B0(N843), .Y(N506) );
  OAI22X1TF U752 ( .A0(N496), .A1(N782), .B0(N199), .B1(N4920), .Y(N501) );
  INVX2TF U753 ( .A(N886), .Y(N4830) );
  AOI21X1TF U754 ( .A0(N427), .A1(REG_A[2]), .B0(N4780), .Y(N886) );
  OAI22X1TF U755 ( .A0(N255), .A1(N222), .B0(N869), .B1(N208), .Y(N4780) );
  NOR4X1TF U756 ( .A(N755), .B(N873), .C(N469), .D(N840), .Y(N877) );
  NOR2X1TF U757 ( .A(N869), .B(N209), .Y(N840) );
  INVX2TF U758 ( .A(N5190), .Y(N869) );
  NOR2X1TF U759 ( .A(N255), .B(N237), .Y(N469) );
  NOR2X1TF U760 ( .A(N785), .B(N219), .Y(N873) );
  NOR2X1TF U761 ( .A(N240), .B(N137), .Y(N755) );
  AOI32X1TF U762 ( .A0(N422), .A1(REG_A[14]), .A2(N199), .B0(N5140), .B1(
        REG_A[14]), .Y(N5110) );
  INVX2TF U763 ( .A(N430), .Y(N285) );
  INVX2TF U764 ( .A(N391), .Y(N388) );
  OAI21X1TF U765 ( .A0(N305), .A1(N229), .B0(N304), .Y(N306) );
  AOI211X1TF U766 ( .A0(N303), .A1(N771), .B0(N302), .C0(N301), .Y(N304) );
  AOI21X1TF U767 ( .A0(N300), .A1(N299), .B0(N843), .Y(N301) );
  AOI22X1TF U768 ( .A0(REG_A[14]), .A1(N5190), .B0(REG_A[13]), .B1(N144), .Y(
        N300) );
  NOR2X1TF U769 ( .A(N298), .B(N782), .Y(N302) );
  INVX2TF U770 ( .A(N420), .Y(N782) );
  NOR2X1TF U771 ( .A(N188), .B(N133), .Y(N861) );
  OAI211X1TF U772 ( .A0(N219), .A1(N138), .B0(N784), .C0(N5180), .Y(N763) );
  NOR2X2TF U773 ( .A(N40), .B(N188), .Y(N863) );
  INVX2TF U774 ( .A(N772), .Y(N339) );
  NOR4BX1TF U775 ( .AN(N776), .B(N766), .C(N5230), .D(N5210), .Y(N772) );
  NOR2X1TF U776 ( .A(N255), .B(N209), .Y(N5210) );
  NOR2X1TF U777 ( .A(N785), .B(N237), .Y(N5230) );
  INVX2TF U778 ( .A(N758), .Y(N785) );
  NOR2X1TF U779 ( .A(N138), .B(N224), .Y(N766) );
  NOR2X2TF U780 ( .A(N38), .B(REG_B[1]), .Y(N5190) );
  NOR2X1TF U781 ( .A(N138), .B(N231), .Y(N5170) );
  NOR2X1TF U782 ( .A(N220), .B(N255), .Y(N765) );
  INVX2TF U783 ( .A(N878), .Y(N303) );
  NAND2X2TF U784 ( .A(N420), .B(N867), .Y(N878) );
  NOR2X2TF U785 ( .A(REG_B[3]), .B(N133), .Y(N867) );
  AOI21X1TF U786 ( .A0(N200), .A1(N259), .B0(N297), .Y(N305) );
  INVX2TF U787 ( .A(N327), .Y(N297) );
  INVX2TF U788 ( .A(N870), .Y(N848) );
  INVX2TF U789 ( .A(N843), .Y(N351) );
  OR2X2TF U790 ( .A(N342), .B(N40), .Y(N843) );
  AND2X2TF U791 ( .A(N1044), .B(N263), .Y(N420) );
  AND2X2TF U792 ( .A(N151), .B(N1014), .Y(N263) );
  INVX2TF U793 ( .A(N889), .Y(N1042) );
  OAI211X1TF U794 ( .A0(N895), .A1(N1043), .B0(N883), .C0(N430), .Y(N541) );
  INVX2TF U795 ( .A(N1044), .Y(N892) );
  NOR3X1TF U796 ( .A(N218), .B(N894), .C(N1017), .Y(N1027) );
  INVX2TF U797 ( .A(N1018), .Y(N894) );
  OR2X2TF U798 ( .A(N267), .B(N266), .Y(N879) );
  NOR2X1TF U799 ( .A(N752), .B(N1043), .Y(N266) );
  INVX2TF U800 ( .A(N425), .Y(N1043) );
  OR2X2TF U801 ( .A(N1021), .B(N39), .Y(N752) );
  AOI21X1TF U802 ( .A0(N265), .A1(N891), .B0(N1016), .Y(N267) );
  INVX2TF U803 ( .A(N1017), .Y(N264) );
  NAND2BX2TF U804 ( .AN(CODE_TYPE[4]), .B(CODE_TYPE[3]), .Y(N1016) );
  AOI211X1TF U805 ( .A0(CODE_TYPE[2]), .A1(N271), .B0(CODE_TYPE[3]), .C0(N270), 
        .Y(N272) );
  INVX2TF U806 ( .A(N1019), .Y(N270) );
  OAI21X1TF U807 ( .A0(N39), .A1(N228), .B0(N268), .Y(N269) );
  INVX2TF U808 ( .A(N549), .Y(N268) );
  NOR2X1TF U809 ( .A(N572), .B(N258), .Y(N549) );
  INVX2TF U810 ( .A(N560), .Y(N261) );
  OAI22X1TF U811 ( .A0(N652), .A1(N154), .B0(N153), .B1(N620), .Y(N1165) );
  OAI22X1TF U812 ( .A0(N668), .A1(N147), .B0(N146), .B1(N231), .Y(N1166) );
  OAI22X1TF U813 ( .A0(N655), .A1(N154), .B0(N153), .B1(N623), .Y(N1060) );
  OAI22X1TF U814 ( .A0(N671), .A1(N147), .B0(N146), .B1(N239), .Y(N1061) );
  OAI22X1TF U815 ( .A0(N660), .A1(N155), .B0(N153), .B1(N628), .Y(N1104) );
  OAI22X1TF U816 ( .A0(N676), .A1(N148), .B0(N146), .B1(N219), .Y(N1105) );
  OAI22X1TF U817 ( .A0(N654), .A1(N155), .B0(N152), .B1(N6220), .Y(N1084) );
  OAI22X1TF U818 ( .A0(N670), .A1(N148), .B0(N145), .B1(N220), .Y(N1085) );
  OAI22X1TF U819 ( .A0(N649), .A1(N155), .B0(N153), .B1(N617), .Y(N1112) );
  OAI22X1TF U820 ( .A0(N665), .A1(N148), .B0(N146), .B1(N210), .Y(N1113) );
  OAI22X1TF U821 ( .A0(N656), .A1(N155), .B0(N153), .B1(N624), .Y(N1176) );
  OAI22X1TF U822 ( .A0(N672), .A1(N148), .B0(N146), .B1(N224), .Y(N1177) );
  OAI22X1TF U823 ( .A0(N648), .A1(N154), .B0(N153), .B1(N616), .Y(N1132) );
  OAI22X1TF U824 ( .A0(N664), .A1(N147), .B0(N145), .B1(N229), .Y(N1133) );
  OAI22X1TF U825 ( .A0(N651), .A1(N154), .B0(N152), .B1(N619), .Y(N1154) );
  OAI22X1TF U826 ( .A0(N667), .A1(N148), .B0(N145), .B1(N227), .Y(N1155) );
  OAI22X1TF U827 ( .A0(N650), .A1(N154), .B0(N153), .B1(N618), .Y(N1078) );
  OAI22X1TF U828 ( .A0(N666), .A1(N148), .B0(N146), .B1(N226), .Y(N1079) );
  OAI22X1TF U829 ( .A0(N661), .A1(N154), .B0(N152), .B1(N629), .Y(N1070) );
  OAI22X1TF U830 ( .A0(N677), .A1(N148), .B0(N145), .B1(N225), .Y(N1071) );
  OAI22X1TF U831 ( .A0(N662), .A1(N154), .B0(N152), .B1(N630), .Y(N1122) );
  OAI22X1TF U832 ( .A0(N678), .A1(N147), .B0(N145), .B1(N208), .Y(N1123) );
  OAI22X1TF U833 ( .A0(N653), .A1(N155), .B0(N152), .B1(N621), .Y(N1094) );
  OAI22X1TF U834 ( .A0(N669), .A1(N148), .B0(N145), .B1(N223), .Y(N1095) );
  OAI22X1TF U835 ( .A0(N663), .A1(N154), .B0(N153), .B1(N631), .Y(N1143) );
  OAI22X1TF U836 ( .A0(N679), .A1(N147), .B0(N146), .B1(N222), .Y(N1144) );
  OAI22X1TF U837 ( .A0(N658), .A1(N155), .B0(N152), .B1(N626), .Y(N1036) );
  OAI22X1TF U838 ( .A0(N657), .A1(N155), .B0(N152), .B1(N625), .Y(N1047) );
  OAI22X1TF U839 ( .A0(N659), .A1(N155), .B0(N152), .B1(N627), .Y(N1053) );
  INVX2TF U840 ( .A(N593), .Y(N5940) );
  AOI21X1TF U841 ( .A0(N259), .A1(N193), .B0(N136), .Y(N357) );
  AOI21X1TF U842 ( .A0(N149), .A1(N831), .B0(N193), .Y(N834) );
  AOI21X1TF U843 ( .A0(N149), .A1(N822), .B0(N194), .Y(N825) );
  AOI21X1TF U844 ( .A0(N150), .A1(N842), .B0(N189), .Y(N847) );
  OAI31X1TF U845 ( .A0(N133), .A1(N875), .A2(N810), .B0(N150), .Y(N811) );
  AOI21X1TF U846 ( .A0(N260), .A1(N190), .B0(N136), .Y(N850) );
  AOI21X1TF U847 ( .A0(N150), .A1(N333), .B0(N190), .Y(N338) );
  AOI22X1TF U848 ( .A0(N168), .A1(REG_A[5]), .B0(N259), .B1(N209), .Y(N333) );
  AOI21X1TF U849 ( .A0(N150), .A1(N757), .B0(N191), .Y(N761) );
  AOI21X1TF U850 ( .A0(N259), .A1(N191), .B0(N136), .Y(N324) );
  AOI21X1TF U851 ( .A0(N427), .A1(N870), .B0(N136), .Y(N809) );
  AOI22X1TF U852 ( .A0(N758), .A1(REG_A[13]), .B0(N143), .B1(REG_A[12]), .Y(
        N759) );
  AOI21X1TF U853 ( .A0(N260), .A1(N195), .B0(N136), .Y(N884) );
  AOI21X1TF U854 ( .A0(N149), .A1(N309), .B0(N195), .Y(N311) );
  AOI22X1TF U855 ( .A0(N424), .A1(REG_A[10]), .B0(N259), .B1(N223), .Y(N309)
         );
  AOI22X1TF U856 ( .A0(N758), .A1(REG_A[15]), .B0(N144), .B1(REG_A[14]), .Y(
        N432) );
  AOI221X1TF U857 ( .A0(N168), .A1(REG_A[12]), .B0(N422), .B1(N227), .C0(N858), 
        .Y(N452) );
  AOI21X1TF U858 ( .A0(N150), .A1(N275), .B0(N198), .Y(N281) );
  AOI22X1TF U859 ( .A0(N168), .A1(REG_A[13]), .B0(N259), .B1(N226), .Y(N275)
         );
  AOI221X1TF U860 ( .A0(N168), .A1(REG_A[14]), .B0(N422), .B1(N210), .C0(N858), 
        .Y(N4920) );
  AOI22X1TF U861 ( .A0(N758), .A1(REG_A[0]), .B0(N143), .B1(REG_A[1]), .Y(
        N5180) );
  AOI21X1TF U862 ( .A0(N150), .A1(N296), .B0(N200), .Y(N307) );
  MXI2X1TF U863 ( .A(N388), .B(N244), .S0(N1195), .Y(N437) );
  OAI32XLTF U864 ( .A0(ZF), .A1(N218), .A2(N891), .B0(N752), .B1(N246), .Y(
        N547) );
  INVX2TF U865 ( .A(N1028), .Y(N596) );
  OAI2BB1X1TF U866 ( .A0N(N186), .A1N(IO_DATAINA[4]), .B0(N379), .Y(N457) );
  OAI2BB1X1TF U867 ( .A0N(N1181), .A1N(N376), .B0(N375), .Y(N377) );
  OAI2BB1X1TF U868 ( .A0N(N186), .A1N(IO_DATAINA[8]), .B0(N382), .Y(N461) );
  NAND2X1TF U869 ( .A(N383), .B(N1183), .Y(N384) );
  OAI2BB1X1TF U870 ( .A0N(N879), .A1N(N519), .B0(N319), .Y(N320) );
  AO21X1TF U871 ( .A0(N259), .A1(N194), .B0(N136), .Y(N318) );
  NAND4X1TF U872 ( .A(N355), .B(N354), .C(N353), .D(N352), .Y(N356) );
  NAND2BX1TF U873 ( .AN(N860), .B(N870), .Y(N352) );
  NAND2BX1TF U874 ( .AN(N844), .B(N351), .Y(N353) );
  AOI2BB1X1TF U875 ( .A0N(N846), .A1N(N845), .B0(N350), .Y(N354) );
  NAND2BX1TF U876 ( .AN(N849), .B(N349), .Y(N350) );
  NAND2X1TF U877 ( .A(N348), .B(REG_A[4]), .Y(N355) );
  AO21X1TF U878 ( .A0(N422), .A1(N189), .B0(N136), .Y(N348) );
  OAI2BB1X1TF U879 ( .A0N(N186), .A1N(IO_DATAINA[7]), .B0(N408), .Y(N5150) );
  AOI2BB1X1TF U880 ( .A0N(N845), .A1N(N807), .B0(N366), .Y(N367) );
  OAI2BB2XLTF U881 ( .B0(N805), .B1(N848), .A0N(N479), .A1N(N253), .Y(N364) );
  OAI2BB1X1TF U882 ( .A0N(N186), .A1N(IO_DATAINA[6]), .B0(N374), .Y(N453) );
  OAI2BB1X1TF U883 ( .A0N(N515), .A1N(N879), .B0(N336), .Y(N337) );
  AO22X1TF U884 ( .A0(N853), .A1(N854), .B0(N870), .B1(N857), .Y(N334) );
  NAND2X1TF U885 ( .A(N516), .B(N879), .Y(N323) );
  AO22X1TF U886 ( .A0(N253), .A1(N478), .B0(N801), .B1(N854), .Y(N340) );
  OAI2BB1X1TF U887 ( .A0N(REG_B[1]), .A1N(N789), .B0(N347), .Y(N371) );
  AOI2BB1X1TF U888 ( .A0N(N787), .A1N(N875), .B0(N346), .Y(N347) );
  NAND3BX1TF U889 ( .AN(N788), .B(N345), .C(N344), .Y(N346) );
  NAND2X1TF U890 ( .A(N252), .B(N511), .Y(N344) );
  OAI2BB2XLTF U891 ( .B0(N342), .B1(N238), .A0N(N870), .A1N(N786), .Y(N343) );
  NAND4X1TF U892 ( .A(N299), .B(N777), .C(N778), .D(N779), .Y(N853) );
  NAND2X1TF U893 ( .A(N1149), .B(IO_STATUS[0]), .Y(N392) );
  OA21XLTF U894 ( .A0(N858), .A1(N328), .B0(REG_B[0]), .Y(N331) );
  OAI2BB2XLTF U895 ( .B0(N882), .B1(N881), .A0N(N888), .A1N(N351), .Y(N310) );
  NAND2X1TF U896 ( .A(N520), .B(N252), .Y(N313) );
  AO22X1TF U897 ( .A0(N351), .A1(N431), .B0(N870), .B1(N862), .Y(N286) );
  AOI222XLTF U898 ( .A0(N448), .A1(N867), .B0(N861), .B1(N832), .C0(N434), 
        .C1(N863), .Y(N456) );
  AO21X1TF U899 ( .A0(N260), .A1(N197), .B0(N5140), .Y(N288) );
  NAND2X1TF U900 ( .A(N522), .B(N252), .Y(N290) );
  OAI2BB1X1TF U901 ( .A0N(N252), .A1N(N523), .B0(N283), .Y(N284) );
  NAND2X1TF U902 ( .A(N420), .B(REG_B[3]), .Y(N821) );
  AO21X1TF U903 ( .A0(N259), .A1(N198), .B0(N5140), .Y(N282) );
  OAI2BB1X1TF U904 ( .A0N(N879), .A1N(N524), .B0(N293), .Y(N294) );
  NAND2X1TF U905 ( .A(N758), .B(REG_A[12]), .Y(N299) );
  MXI2X1TF U906 ( .A(N259), .B(N168), .S0(REG_A[15]), .Y(N296) );
  NAND2X1TF U907 ( .A(N1044), .B(N39), .Y(N265) );
  NAND2BX1TF U908 ( .AN(N272), .B(N542), .Y(N273) );
  AOI2BB1X1TF U909 ( .A0N(N1044), .A1N(N269), .B0(N212), .Y(N274) );
  OAI2BB1X1TF U910 ( .A0N(N212), .A1N(N572), .B0(N261), .Y(N262) );
  CLKBUFX2TF U911 ( .A(N409), .Y(N254) );
  CLKBUFX2TF U912 ( .A(N1189), .Y(N257) );
  CLKBUFX2TF U913 ( .A(N1186), .Y(N256) );
  NAND2X1TF U914 ( .A(N5190), .B(REG_A[12]), .Y(N768) );
  NAND2X1TF U915 ( .A(N758), .B(REG_A[10]), .Y(N767) );
  OAI221XLTF U916 ( .A0(N38), .A1(REG_A[0]), .B0(REG_B[0]), .B1(REG_A[1]), 
        .C0(N187), .Y(N781) );
  NAND2X1TF U917 ( .A(N427), .B(REG_A[9]), .Y(N778) );
  NAND2X1TF U918 ( .A(CODE_TYPE[4]), .B(N562), .Y(N1019) );
  NAND2X1TF U919 ( .A(N5190), .B(REG_A[11]), .Y(N760) );
  NAND2X1TF U920 ( .A(N5190), .B(REG_A[13]), .Y(N460) );
  OAI222X1TF U921 ( .A0(N141), .A1(N419), .B0(N140), .B1(N417), .C0(N423), 
        .C1(N251), .Y(N470) );
  NAND2X1TF U922 ( .A(N144), .B(REG_A[12]), .Y(N465) );
  NAND2X1TF U923 ( .A(N758), .B(REG_A[11]), .Y(N827) );
  NAND2X1TF U924 ( .A(N794), .B(N133), .Y(N753) );
  NAND2X1TF U925 ( .A(N427), .B(REG_A[10]), .Y(N473) );
  NAND2X1TF U926 ( .A(REG_A[9]), .B(N5190), .Y(N829) );
  NAND2X1TF U927 ( .A(N758), .B(REG_A[7]), .Y(N841) );
  NAND4X1TF U928 ( .A(N756), .B(N473), .C(N829), .D(N841), .Y(N888) );
  AOI222XLTF U929 ( .A0(N4870), .A1(N863), .B0(N888), .B1(N867), .C0(N4830), 
        .C1(N861), .Y(N496) );
  OAI222X1TF U930 ( .A0(N140), .A1(N419), .B0(N142), .B1(N415), .C0(N418), 
        .C1(N251), .Y(N4880) );
  NAND2X1TF U931 ( .A(N758), .B(REG_A[8]), .Y(N775) );
  NAND2X1TF U932 ( .A(N5190), .B(REG_A[10]), .Y(N779) );
  NAND4BBX1TF U933 ( .AN(N765), .BN(N5170), .C(N775), .D(N779), .Y(N771) );
  NAND2X1TF U934 ( .A(N5190), .B(REG_A[2]), .Y(N784) );
  NAND2X1TF U935 ( .A(REG_A[6]), .B(N5190), .Y(N776) );
  NAND3X1TF U936 ( .A(N215), .B(N221), .C(N211), .Y(N540) );
  NAND2X1TF U937 ( .A(N743), .B(START), .Y(N741) );
  NOR4XLTF U938 ( .A(N258), .B(N1021), .C(N890), .D(N564), .Y(N173) );
  NAND2X1TF U939 ( .A(N716), .B(I_ADDR[4]), .Y(N717) );
  NAND2X1TF U940 ( .A(N721), .B(I_ADDR[6]), .Y(N726) );
  NOR2BX1TF U941 ( .AN(N738), .B(N737), .Y(N174) );
  NAND2X1TF U942 ( .A(N232), .B(N215), .Y(N544) );
  NOR4XLTF U943 ( .A(N752), .B(N544), .C(N221), .D(N890), .Y(N622) );
  NAND2X1TF U944 ( .A(N39), .B(N572), .Y(N751) );
  NOR2BX1TF U945 ( .AN(N551), .B(N737), .Y(N550) );
  NAND2X1TF U946 ( .A(N566), .B(N551), .Y(N724) );
  AO22X1TF U947 ( .A0(D_ADDR[8]), .A1(N729), .B0(I_ADDR[8]), .B1(N722), .Y(
        N553) );
  NAND2X1TF U948 ( .A(N730), .B(N731), .Y(N555) );
  OAI221XLTF U949 ( .A0(N39), .A1(N212), .B0(N258), .B1(N425), .C0(N572), .Y(
        N556) );
  NAND2X1TF U950 ( .A(I_ADDR[1]), .B(I_ADDR[2]), .Y(N713) );
  NAND3X1TF U951 ( .A(N730), .B(N232), .C(N215), .Y(N739) );
  NOR4XLTF U952 ( .A(N558), .B(IO_STATUS[0]), .C(IO_STATUS[1]), .D(N733), .Y(
        N736) );
  NAND2X1TF U954 ( .A(N243), .B(N747), .Y(N1030) );
  NAND2X1TF U955 ( .A(N212), .B(N1044), .Y(N1015) );
  NAND2X1TF U956 ( .A(N880), .B(REG_B[3]), .Y(N795) );
  NAND2X1TF U957 ( .A(N427), .B(REG_A[15]), .Y(N810) );
  NAND2X1TF U958 ( .A(N880), .B(N863), .Y(N851) );
  NAND2X1TF U959 ( .A(N420), .B(N863), .Y(N885) );
  NAND4X1TF U960 ( .A(N776), .B(N775), .C(N774), .D(N773), .Y(N857) );
  AOI222XLTF U961 ( .A0(N857), .A1(N867), .B0(N853), .B1(N863), .C0(N780), 
        .C1(N861), .Y(N787) );
  NAND2X1TF U962 ( .A(N144), .B(REG_A[3]), .Y(N783) );
  AOI2BB2X1TF U963 ( .B0(REG_A[3]), .B1(N818), .A0N(N188), .A1N(N817), .Y(N819) );
  NAND4BX1TF U964 ( .AN(N830), .B(N829), .C(N828), .D(N827), .Y(N866) );
  AOI222XLTF U965 ( .A0(N868), .A1(N867), .B0(N866), .B1(N863), .C0(N862), 
        .C1(N861), .Y(N876) );
  NAND2X1TF U966 ( .A(N188), .B(N880), .Y(N882) );
  NAND2X1TF U967 ( .A(N1024), .B(N919), .Y(N1185) );
  AOI2BB2X1TF U968 ( .B0(IO_DATAINA[2]), .B1(N186), .A0N(N411), .A1N(N142), 
        .Y(N1076) );
  NAND3X1TF U969 ( .A(N1131), .B(N1130), .C(N1129), .Y(N493) );
  AOI2BB2X1TF U970 ( .B0(N406), .B1(N1198), .A0N(N1198), .A1N(I_DATAIN[7]), 
        .Y(N532) );
  OAI2BB2XLTF U971 ( .B0(N166), .B1(N405), .A0N(N166), .A1N(I_DATAIN[6]), .Y(
        N533) );
  OAI2BB2XLTF U972 ( .B0(N166), .B1(N404), .A0N(N166), .A1N(I_DATAIN[5]), .Y(
        N534) );
  AO22X1TF U973 ( .A0(N1198), .A1(N236), .B0(N166), .B1(I_DATAIN[4]), .Y(N535)
         );
  AOI2BB2X1TF U974 ( .B0(N402), .B1(N1198), .A0N(N1198), .A1N(I_DATAIN[3]), 
        .Y(N536) );
  OAI2BB2XLTF U975 ( .B0(N165), .B1(N213), .A0N(N166), .A1N(I_DATAIN[2]), .Y(
        N537) );
  OAI2BB2XLTF U976 ( .B0(N165), .B1(N217), .A0N(N166), .A1N(I_DATAIN[1]), .Y(
        N538) );
  OAI2BB2XLTF U977 ( .B0(N165), .B1(N235), .A0N(N166), .A1N(I_DATAIN[0]), .Y(
        N539) );
endmodule


module SCPU_SRAM_8BIT_ALU_SPI_TOP_VG ( CLK, RST_N, CTRL_MODE, CTRL_BGN, CPU_BGN, 
        LOAD_N, CTRL_SI, ADC_PI, CTRL_RDY, CTRL_SO, NXT, SCLK1, SCLK2, LAT, 
        SPI_SO );
  input [1:0] CTRL_MODE;
  input [9:0] ADC_PI;
  output [1:0] NXT;
  input CLK, RST_N, CTRL_BGN, CPU_BGN, LOAD_N, CTRL_SI;
  output CTRL_RDY, CTRL_SO, SCLK1, SCLK2, LAT, SPI_SO;
  wire   CEN_AFTER_MUX, WEN_AFTER_MUX, I_CLK, I_RST_N, I_CTRL_BGN, I_CPU_BGN,
         I_LOAD_N, I_CTRL_SI, I_CTRL_SO, I_SCLK1, I_SCLK2, I_SPI_SO,
         SCPU_CTRL_SPI_CEN, \SCPU_CTRL_SPI_IO_DATAOUTB[0] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[1] , \SCPU_CTRL_SPI_IO_DATAOUTB[2] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[3] , \SCPU_CTRL_SPI_IO_DATAOUTB[4] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[5] , \SCPU_CTRL_SPI_IO_DATAOUTB[6] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[7] , \SCPU_CTRL_SPI_IO_DATAOUTB[8] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[9] , \SCPU_CTRL_SPI_IO_DATAOUTB[10] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[11] , \SCPU_CTRL_SPI_IO_DATAOUTB[12] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[0] , \SCPU_CTRL_SPI_IO_DATAOUTA[1] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[2] , \SCPU_CTRL_SPI_IO_DATAOUTA[3] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[4] , \SCPU_CTRL_SPI_IO_DATAOUTA[5] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[6] , \SCPU_CTRL_SPI_IO_DATAOUTA[7] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[8] , \SCPU_CTRL_SPI_IO_DATAOUTA[9] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[10] , \SCPU_CTRL_SPI_IO_DATAOUTA[11] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[12] , \SCPU_CTRL_SPI_IO_CONTROL[0] ,
         \SCPU_CTRL_SPI_IO_CONTROL[1] , \SCPU_CTRL_SPI_IO_CONTROL[2] ,
         \SCPU_CTRL_SPI_IO_CONTROL[3] , \SCPU_CTRL_SPI_IO_CONTROL[4] ,
         \SCPU_CTRL_SPI_IO_CONTROL[5] , \SCPU_CTRL_SPI_IO_CONTROL[6] ,
         SCPU_CTRL_SPI_D_WE, SCPU_CTRL_SPI_IS_I_ADDR, SCPU_CTRL_SPI_CCT_N57,
         SCPU_CTRL_SPI_CCT_N56, SCPU_CTRL_SPI_CCT_N55, SCPU_CTRL_SPI_CCT_N53,
         SCPU_CTRL_SPI_CCT_N52, SCPU_CTRL_SPI_CCT_N51,
         SCPU_CTRL_SPI_CCT_IS_SHIFT, \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[3] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[5] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[7] , \SCPU_CTRL_SPI_CCT_REG_BITS[1] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[2] , \SCPU_CTRL_SPI_CCT_REG_BITS[3] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[4] , \SCPU_CTRL_SPI_CCT_REG_BITS[5] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[6] , \SCPU_CTRL_SPI_CCT_REG_BITS[7] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[8] , \SCPU_CTRL_SPI_CCT_REG_BITS[9] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[10] , \SCPU_CTRL_SPI_CCT_REG_BITS[11] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[12] , \SCPU_CTRL_SPI_CCT_REG_BITS[13] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[14] , \SCPU_CTRL_SPI_CCT_REG_BITS[15] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[16] , \SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ,
         SCPU_CTRL_SPI_PUT_N110, SCPU_CTRL_SPI_PUT_N109,
         SCPU_CTRL_SPI_PUT_N108, \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] , SCPU_CTRL_SPI_PUT_N27,
         SCPU_CTRL_SPI_PUT_IS_ADDR_LEN_NZ, \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ,
         \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ,
         \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] ,
         \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[4] , \SCPU_CTRL_SPI_PUT_SPI_STATE[0] ,
         \SCPU_CTRL_SPI_PUT_SPI_STATE[1] , \SCPU_CTRL_SPI_PUT_CNT_STATE[0] ,
         \SCPU_CTRL_SPI_PUT_CNT_STATE[1] , \SCPU_CTRL_SPI_PUT_CNT_STATE[2] ,
         N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45,
         N46, N81, N82, N83, N84, N85, N86, N87, N88, N89, N93, N95, N103,
         N105, N161, N167, N168, N192, N193, N194, N195, N196, N197, N198,
         N199, N200, N201, N202, N203, N204, N205, N206, N207, N208, N209,
         N210, N211, N212, N213, N215, N216, N217, N218, N219, N221, N222,
         N223, N224, N225, N236, N237, N238, N263, N264, N265, N266, N267,
         N268, N271, N272, N273, N274, N275, N276, N277, N278, N279, N280,
         N281, N282, N283, N284, N285, N286, N287, N288, N289, N290, N291,
         N292, N293, N294, N295, N296, N297, N298, N299, N300, N301, N302,
         N303, N304, N305, N306, N307, N308, N309, N310, N311, N312, N313,
         N314, N315, N316, N317, N318, N319, N320, N321, N322, N323, N324,
         N325, N326, N327, N328, N329, N330, N331, N332, N333, N334, N335,
         N336, N337, N338, N339, N340, N341, N342, N343, N344, N345, N346,
         N347, N348, N349, N350, N351, N352, N353, N354, N355, N356, N357,
         N358, N359, N360, N361, N362, N363, N364, N365, N366, N367, N368,
         N369, N370, N371, N372, N373, N374, N375, N376, N377, N378, N379,
         N380, N381, N382, N383, N384, N385, N386, N387, N388, N389, N390,
         N391, N392, N393, N394, N395, N396, N397, N398, N399, N400, N401,
         N402, N403, N404, N405, N406, N407, N408, N409, N410, N411, N412,
         N413, N414, N415, N416, N417, N418, N419, N420, N421, N422, N423,
         N424;
  wire   [8:0] A_AFTER_MUX;
  wire   [7:0] D_AFTER_MUX;
  wire   [7:0] Q_FROM_SRAM;
  wire   [1:0] I_CTRL_MODE;
  wire   [9:0] I_ADC_PI;
  wire   [1:0] I_NXT;
  wire   [8:0] SCPU_CTRL_SPI_A_SPI;
  wire   [12:0] SCPU_CTRL_SPI_POUT;
  wire   [12:0] SCPU_CTRL_SPI_FOUT;
  wire   [9:0] SCPU_CTRL_SPI_IO_OFFSET;
  wire   [12:0] SCPU_CTRL_SPI_IO_DATAINA;
  wire   [0:0] SCPU_CTRL_SPI_IO_STATUS;
  wire   [7:0] SCPU_CTRL_SPI_D_DATAOUT;
  wire   [8:1] SCPU_CTRL_SPI_D_ADDR;
  wire   [8:0] SCPU_CTRL_SPI_I_ADDR;
  wire   [7:0] SCPU_CTRL_SPI_D_DATAIN;
  wire   [7:0] SCPU_CTRL_SPI_I_DATAIN;
  wire   [7:1] SCPU_CTRL_SPI_PUT_SRAM_REGS;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21;

  RA1SHD_IBM512X8 sram ( .Q(Q_FROM_SRAM), .A(A_AFTER_MUX), .D(D_AFTER_MUX), 
        .CLK(I_CLK), .CEN(CEN_AFTER_MUX), .WEN(WEN_AFTER_MUX) );
  PIC ipad_clk ( .IE(1'b1), .P(CLK), .Y(I_CLK) );
  PIC ipad_rst_n ( .IE(1'b1), .P(RST_N), .Y(I_RST_N) );
  PIC ipad_ctrl_mode0 ( .IE(1'b1), .P(CTRL_MODE[0]), .Y(I_CTRL_MODE[0]) );
  PIC ipad_ctrl_mode1 ( .IE(1'b1), .P(CTRL_MODE[1]), .Y(I_CTRL_MODE[1]) );
  PIC ipad_ctrl_bgn ( .IE(1'b1), .P(CTRL_BGN), .Y(I_CTRL_BGN) );
  PIC ipad_cpu_str ( .IE(1'b1), .P(CPU_BGN), .Y(I_CPU_BGN) );
  PIC ipad_load_n ( .IE(1'b1), .P(LOAD_N), .Y(I_LOAD_N) );
  PIC ipad_ctrl_si ( .IE(1'b1), .P(CTRL_SI), .Y(I_CTRL_SI) );
  PIC ipad_adc_pi0 ( .IE(1'b1), .P(ADC_PI[0]), .Y(I_ADC_PI[0]) );
  PIC ipad_adc_pi1 ( .IE(1'b1), .P(ADC_PI[1]), .Y(I_ADC_PI[1]) );
  PIC ipad_adc_pi2 ( .IE(1'b1), .P(ADC_PI[2]), .Y(I_ADC_PI[2]) );
  PIC ipad_adc_pi3 ( .IE(1'b1), .P(ADC_PI[3]), .Y(I_ADC_PI[3]) );
  PIC ipad_adc_pi4 ( .IE(1'b1), .P(ADC_PI[4]), .Y(I_ADC_PI[4]) );
  PIC ipad_adc_pi5 ( .IE(1'b1), .P(ADC_PI[5]), .Y(I_ADC_PI[5]) );
  PIC ipad_adc_pi6 ( .IE(1'b1), .P(ADC_PI[6]), .Y(I_ADC_PI[6]) );
  PIC ipad_adc_pi7 ( .IE(1'b1), .P(ADC_PI[7]), .Y(I_ADC_PI[7]) );
  PIC ipad_adc_pi8 ( .IE(1'b1), .P(ADC_PI[8]), .Y(I_ADC_PI[8]) );
  PIC ipad_adc_pi9 ( .IE(1'b1), .P(ADC_PI[9]), .Y(I_ADC_PI[9]) );
  POC8B opad_ctrl_rdy ( .A(N223), .P(CTRL_RDY) );
  POC8B opad_ctrl_so ( .A(I_CTRL_SO), .P(CTRL_SO) );
  POC8B opad_nxt0 ( .A(I_NXT[0]), .P(NXT[0]) );
  POC8B opad_nxt1 ( .A(I_NXT[1]), .P(NXT[1]) );
  POC8B opad_sclk1 ( .A(I_SCLK1), .P(SCLK1) );
  POC8B opad_sclk2 ( .A(I_SCLK2), .P(SCLK2) );
  POC8B opad_lat ( .A(N225), .P(LAT) );
  POC8B opad_spi_so ( .A(I_SPI_SO), .P(SPI_SO) );
  SHARE_SUPERALU_VG \scpu_ctrl_spi/ALU_01  ( .CLK(I_CLK), .RST_N(I_RST_N), .X_IN(
        {\SCPU_CTRL_SPI_IO_DATAOUTA[12] , \SCPU_CTRL_SPI_IO_DATAOUTA[11] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[10] , \SCPU_CTRL_SPI_IO_DATAOUTA[9] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[8] , \SCPU_CTRL_SPI_IO_DATAOUTA[7] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[6] , \SCPU_CTRL_SPI_IO_DATAOUTA[5] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[4] , \SCPU_CTRL_SPI_IO_DATAOUTA[3] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[2] , \SCPU_CTRL_SPI_IO_DATAOUTA[1] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[0] }), .Y_IN({
        \SCPU_CTRL_SPI_IO_DATAOUTB[12] , \SCPU_CTRL_SPI_IO_DATAOUTB[11] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[10] , \SCPU_CTRL_SPI_IO_DATAOUTB[9] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[8] , \SCPU_CTRL_SPI_IO_DATAOUTB[7] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[6] , \SCPU_CTRL_SPI_IO_DATAOUTB[5] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[4] , \SCPU_CTRL_SPI_IO_DATAOUTB[3] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[2] , \SCPU_CTRL_SPI_IO_DATAOUTB[1] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[0] }), .ALU_START(N265), .ALU_TYPE({
        \SCPU_CTRL_SPI_IO_CONTROL[4] , \SCPU_CTRL_SPI_IO_CONTROL[3] , 
        \SCPU_CTRL_SPI_IO_CONTROL[2] }), .MODE_TYPE({
        \SCPU_CTRL_SPI_IO_CONTROL[1] , \SCPU_CTRL_SPI_IO_CONTROL[0] }), 
        .OFFSET(SCPU_CTRL_SPI_IO_OFFSET), .FOUT(SCPU_CTRL_SPI_FOUT), .POUT(
        SCPU_CTRL_SPI_POUT), .ALU_IS_DONE(SCPU_CTRL_SPI_IO_STATUS[0]) );
  SERIAL_CPU_8BIT_VG \scpu_ctrl_spi/uut  ( .CLK(I_CLK), .ENABLE(1'b0), .RST_N(
        I_RST_N), .START(I_CPU_BGN), .I_DATAIN(SCPU_CTRL_SPI_I_DATAIN), 
        .D_DATAIN(SCPU_CTRL_SPI_D_DATAIN), .IS_I_ADDR(SCPU_CTRL_SPI_IS_I_ADDR), 
        .NXT(I_NXT), .I_ADDR(SCPU_CTRL_SPI_I_ADDR), .D_ADDR({
        SCPU_CTRL_SPI_D_ADDR, SYNOPSYS_UNCONNECTED__0}), .D_WE(
        SCPU_CTRL_SPI_D_WE), .D_DATAOUT(SCPU_CTRL_SPI_D_DATAOUT), .IO_STATUS({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, N224, SCPU_CTRL_SPI_IO_STATUS[0]}), .IO_CONTROL({
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, \SCPU_CTRL_SPI_IO_CONTROL[6] , 
        \SCPU_CTRL_SPI_IO_CONTROL[5] , \SCPU_CTRL_SPI_IO_CONTROL[4] , 
        \SCPU_CTRL_SPI_IO_CONTROL[3] , \SCPU_CTRL_SPI_IO_CONTROL[2] , 
        \SCPU_CTRL_SPI_IO_CONTROL[1] , \SCPU_CTRL_SPI_IO_CONTROL[0] }), 
        .IO_DATAINA({1'b0, 1'b0, 1'b0, SCPU_CTRL_SPI_IO_DATAINA}), 
        .IO_DATAINB({1'b0, 1'b0, 1'b0, SCPU_CTRL_SPI_POUT}), .IO_DATAOUTA({
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, \SCPU_CTRL_SPI_IO_DATAOUTA[12] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[11] , \SCPU_CTRL_SPI_IO_DATAOUTA[10] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[9] , \SCPU_CTRL_SPI_IO_DATAOUTA[8] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[7] , \SCPU_CTRL_SPI_IO_DATAOUTA[6] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[5] , \SCPU_CTRL_SPI_IO_DATAOUTA[4] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[3] , \SCPU_CTRL_SPI_IO_DATAOUTA[2] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[1] , \SCPU_CTRL_SPI_IO_DATAOUTA[0] }), 
        .IO_DATAOUTB({SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, \SCPU_CTRL_SPI_IO_DATAOUTB[12] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[11] , \SCPU_CTRL_SPI_IO_DATAOUTB[10] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[9] , \SCPU_CTRL_SPI_IO_DATAOUTB[8] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[7] , \SCPU_CTRL_SPI_IO_DATAOUTB[6] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[5] , \SCPU_CTRL_SPI_IO_DATAOUTB[4] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[3] , \SCPU_CTRL_SPI_IO_DATAOUTB[2] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[1] , \SCPU_CTRL_SPI_IO_DATAOUTB[0] }), 
        .IO_OFFSET({SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SCPU_CTRL_SPI_IO_OFFSET}) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[7]  ( .D(N161), .RN(
        SCPU_CTRL_SPI_CCT_N57), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[7] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[5]  ( .D(N161), .RN(
        SCPU_CTRL_SPI_CCT_N55), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[5] ), .QN(N284) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[3]  ( .D(N161), .RN(
        SCPU_CTRL_SPI_CCT_N53), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[3] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[2]  ( .D(N161), .RN(
        SCPU_CTRL_SPI_CCT_N52), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[1]  ( .D(N161), .RN(
        SCPU_CTRL_SPI_CCT_N51), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[6]  ( .D(N161), .RN(
        SCPU_CTRL_SPI_CCT_N56), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[16]  ( .D(I_CTRL_SI), .E(N267), 
        .CK(I_CLK), .Q(\SCPU_CTRL_SPI_CCT_REG_BITS[16] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[15]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[16] ), .E(N267), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[15] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[14]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[15] ), .E(N267), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[14] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[13]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[14] ), .E(N267), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[13] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[12]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[13] ), .E(N267), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[12] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[11]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[12] ), .E(N267), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[11] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[10]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[11] ), .E(N267), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[10] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[9]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[10] ), .E(N267), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[9] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[8]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[9] ), .E(N267), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[8] ) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[2]  ( .D(N40), .CK(I_CLK), 
        .SN(N39), .RN(N38), .QN(N286) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[4]  ( .D(N46), .CK(I_CLK), 
        .SN(N45), .RN(N44), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[4] ), .QN(N280)
         );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[1]  ( .D(N37), .CK(I_CLK), 
        .SN(N36), .RN(N35), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ), .QN(N277)
         );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[3]  ( .D(N43), .CK(I_CLK), 
        .SN(N42), .RN(N41), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] ), .QN(N274)
         );
  DFFSX2TF \scpu_ctrl_spi/put/cnt_state_reg[0]  ( .D(SCPU_CTRL_SPI_PUT_N108), 
        .CK(I_CLK), .SN(\SCPU_CTRL_SPI_IO_CONTROL[6] ), .Q(
        \SCPU_CTRL_SPI_PUT_CNT_STATE[0] ), .QN(N272) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[7]  ( .D(N192), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[7] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[6]  ( .D(N193), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[6] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[5]  ( .D(N194), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[5] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[4]  ( .D(N195), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[4] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[3]  ( .D(N196), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[3] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[2]  ( .D(N197), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[2] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[1]  ( .D(N198), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[1] ) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[7]  ( .D(N207), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[7]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[6]  ( .D(N201), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[6]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[5]  ( .D(N202), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[5]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[4]  ( .D(N203), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[4]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[3]  ( .D(N204), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[3]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[2]  ( .D(N205), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[2]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[1]  ( .D(N206), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[1]) );
  DFFTRX1TF \scpu_ctrl_spi/cct/is_shift_reg  ( .D(N167), .RN(N168), .CK(I_CLK), 
        .QN(SCPU_CTRL_SPI_CCT_IS_SHIFT) );
  DFFQX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[4]  ( .D(N218), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[0]  ( .D(N217), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[0]  ( .D(N200), .CK(I_CLK), .Q(
        I_SPI_SO) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[0]  ( .D(N199), .CK(I_CLK), .Q(
        I_CTRL_SO) );
  DFFXLTF \scpu_ctrl_spi/cct/ctrl_state_reg[0]  ( .D(N219), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .QN(N288) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[0]  ( .D(N34), .CK(I_CLK), 
        .SN(N33), .RN(N32), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ) );
  DFFNSRX4TF \scpu_ctrl_spi/put/spi_MUX_reg  ( .D(N216), .CKN(I_CLK), .SN(1'b1), .RN(1'b1), .Q(N300), .QN(N105) );
  DFFNSRX1TF \scpu_ctrl_spi/cct/D_WE_reg  ( .D(N221), .CKN(I_CLK), .SN(1'b1), 
        .RN(1'b1), .QN(N281) );
  DFFNSRX1TF \scpu_ctrl_spi/put/sram_addr_reg[5]  ( .D(N86), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[5]), .QN(N276) );
  DFFNSRX1TF \scpu_ctrl_spi/put/sram_addr_reg[6]  ( .D(N87), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[6]), .QN(N282) );
  DFFNSRX1TF \scpu_ctrl_spi/put/sram_addr_reg[7]  ( .D(N88), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[7]), .QN(N283) );
  DFFNSRXLTF \scpu_ctrl_spi/cct/CEN_reg  ( .D(N222), .CKN(I_CLK), .SN(1'b1), 
        .RN(1'b1), .Q(SCPU_CTRL_SPI_CEN) );
  DFFNSRXLTF \scpu_ctrl_spi/put/is_addr_len_nz_reg  ( .D(SCPU_CTRL_SPI_PUT_N27), .CKN(I_CLK), .SN(1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_PUT_IS_ADDR_LEN_NZ) );
  DFFNSRXLTF \scpu_ctrl_spi/put/sram_addr_reg[8]  ( .D(N89), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[8]) );
  EDFFTRXLTF \scpu_ctrl_spi/cct/ctrl_state_reg[1]  ( .RN(I_CTRL_BGN), .D(1'b1), 
        .E(N238), .CK(I_CLK), .Q(N279), .QN(N95) );
  DFFRX1TF \scpu_ctrl_spi/put/cnt_state_reg[2]  ( .D(SCPU_CTRL_SPI_PUT_N110), 
        .CK(I_CLK), .RN(N291), .Q(\SCPU_CTRL_SPI_PUT_CNT_STATE[2] ) );
  DFFRX1TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[1]  ( .D(N209), .CK(I_CLK), 
        .RN(N291), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ) );
  DFFRX1TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[2]  ( .D(N210), .CK(I_CLK), 
        .RN(N291), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ) );
  DFFRX2TF \scpu_ctrl_spi/put/cnt_state_reg[1]  ( .D(SCPU_CTRL_SPI_PUT_N109), 
        .CK(I_CLK), .RN(N291), .Q(\SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .QN(N275)
         );
  DFFRX2TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[0]  ( .D(N208), .CK(I_CLK), 
        .RN(N291), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .QN(N278) );
  DFFRX2TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[3]  ( .D(N211), .CK(I_CLK), 
        .RN(\SCPU_CTRL_SPI_IO_CONTROL[6] ), .Q(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ), .QN(N287) );
  DFFRX2TF \scpu_ctrl_spi/put/spi_state_reg[2]  ( .D(N215), .CK(I_CLK), .RN(
        \SCPU_CTRL_SPI_IO_CONTROL[6] ), .Q(N271), .QN(N103) );
  DFFRX2TF \scpu_ctrl_spi/put/spi_state_reg[1]  ( .D(N213), .CK(I_CLK), .RN(
        \SCPU_CTRL_SPI_IO_CONTROL[6] ), .Q(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), 
        .QN(N289) );
  DFFRX2TF \scpu_ctrl_spi/put/spi_state_reg[0]  ( .D(N212), .CK(I_CLK), .RN(
        \SCPU_CTRL_SPI_IO_CONTROL[6] ), .Q(\SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), 
        .QN(N273) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[1]  ( .D(N82), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[1]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[3]  ( .D(N84), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[3]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[2]  ( .D(N83), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[2]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[4]  ( .D(N85), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[4]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[0]  ( .D(N81), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[0]), .QN(N285) );
  NOR3BX2TF U245 ( .AN(N286), .B(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .C(
        \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ), .Y(N423) );
  CLKBUFX2TF U246 ( .A(N292), .Y(N293) );
  AND2X2TF U247 ( .A(N320), .B(N281), .Y(N321) );
  AND2X1TF U248 ( .A(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .B(SCPU_CTRL_SPI_FOUT[10]), .Y(SCPU_CTRL_SPI_IO_DATAINA[10]) );
  AND2X1TF U249 ( .A(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .B(SCPU_CTRL_SPI_FOUT[11]), .Y(SCPU_CTRL_SPI_IO_DATAINA[11]) );
  AND2X1TF U250 ( .A(N265), .B(SCPU_CTRL_SPI_FOUT[12]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[12]) );
  OAI22X1TF U251 ( .A0(SCPU_CTRL_SPI_PUT_IS_ADDR_LEN_NZ), .A1(N419), .B0(N333), 
        .B1(N271), .Y(N236) );
  AOI21X1TF U252 ( .A0(N333), .A1(N271), .B0(N236), .Y(N237) );
  AOI22X1TF U253 ( .A0(N337), .A1(N237), .B0(N103), .B1(N339), .Y(N215) );
  OA21XLTF U254 ( .A0(N268), .A1(I_CTRL_MODE[0]), .B0(N322), .Y(N238) );
  AND2X1TF U269 ( .A(N418), .B(N291), .Y(SCPU_CTRL_SPI_PUT_N27) );
  NAND3X1TF U270 ( .A(SCPU_CTRL_SPI_CCT_IS_SHIFT), .B(N95), .C(N268), .Y(N93)
         );
  NOR2X4TF U271 ( .A(SCPU_CTRL_SPI_CEN), .B(N263), .Y(N320) );
  NAND2XLTF U272 ( .A(N272), .B(N275), .Y(N386) );
  AOI22X1TF U273 ( .A0(N317), .A1(SCPU_CTRL_SPI_D_ADDR[8]), .B0(N320), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[16] ), .Y(N318) );
  AOI22X1TF U274 ( .A0(N317), .A1(SCPU_CTRL_SPI_D_ADDR[7]), .B0(N320), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[15] ), .Y(N313) );
  AOI22X1TF U275 ( .A0(N317), .A1(SCPU_CTRL_SPI_D_ADDR[6]), .B0(N320), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[14] ), .Y(N311) );
  AOI22X1TF U276 ( .A0(N317), .A1(SCPU_CTRL_SPI_D_ADDR[5]), .B0(N320), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[13] ), .Y(N309) );
  AOI22X1TF U277 ( .A0(N317), .A1(SCPU_CTRL_SPI_D_ADDR[4]), .B0(N320), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[12] ), .Y(N307) );
  AOI22X1TF U278 ( .A0(N317), .A1(SCPU_CTRL_SPI_D_ADDR[3]), .B0(N320), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[11] ), .Y(N305) );
  AOI22X1TF U279 ( .A0(N317), .A1(SCPU_CTRL_SPI_D_ADDR[2]), .B0(N320), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[10] ), .Y(N303) );
  AOI22X1TF U280 ( .A0(N317), .A1(SCPU_CTRL_SPI_D_ADDR[1]), .B0(N320), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[9] ), .Y(N301) );
  NAND2XLTF U281 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[4] ), .B(N294), .Y(N45) );
  NAND2XLTF U282 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[3] ), .B(N294), .Y(N42) );
  NAND2XLTF U283 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[2] ), .B(N294), .Y(N39) );
  NAND2BXLTF U284 ( .AN(\SCPU_CTRL_SPI_IO_DATAOUTB[4] ), .B(N292), .Y(N44) );
  NAND2BXLTF U285 ( .AN(\SCPU_CTRL_SPI_IO_DATAOUTB[3] ), .B(N292), .Y(N41) );
  NAND2BXLTF U286 ( .AN(\SCPU_CTRL_SPI_IO_DATAOUTB[0] ), .B(N292), .Y(N32) );
  OAI211XLTF U287 ( .A0(\SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .A1(N336), .B0(N337), .C0(N271), .Y(N335) );
  INVX1TF U288 ( .A(N323), .Y(N324) );
  NAND2XLTF U289 ( .A(N404), .B(SCPU_CTRL_SPI_A_SPI[3]), .Y(N403) );
  NAND2BXLTF U290 ( .AN(\SCPU_CTRL_SPI_IO_DATAOUTB[2] ), .B(N417), .Y(N38) );
  NAND2XLTF U291 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[1] ), .B(N417), .Y(N36) );
  NAND2BXLTF U292 ( .AN(\SCPU_CTRL_SPI_IO_DATAOUTB[1] ), .B(N417), .Y(N35) );
  NAND2XLTF U293 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[0] ), .B(N417), .Y(N33) );
  NAND2BX2TF U294 ( .AN(SCPU_CTRL_SPI_IS_I_ADDR), .B(N263), .Y(N374) );
  INVX2TF U295 ( .A(I_CTRL_BGN), .Y(N263) );
  INVX2TF U296 ( .A(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .Y(N290) );
  OR2X2TF U297 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ), .B(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .Y(N295) );
  NAND2XLTF U298 ( .A(SCPU_CTRL_SPI_A_SPI[0]), .B(SCPU_CTRL_SPI_A_SPI[1]), .Y(
        N410) );
  CLKBUFX2TF U299 ( .A(\SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .Y(N268) );
  INVX2TF U300 ( .A(I_CTRL_BGN), .Y(N264) );
  INVX2TF U301 ( .A(N290), .Y(N265) );
  INVX2TF U302 ( .A(N93), .Y(N266) );
  INVX2TF U303 ( .A(N93), .Y(N267) );
  NOR3X4TF U304 ( .A(I_CTRL_BGN), .B(N293), .C(N351), .Y(N360) );
  NOR3X1TF U305 ( .A(N268), .B(N279), .C(N264), .Y(N325) );
  NAND4BX2TF U306 ( .AN(N222), .B(I_CTRL_BGN), .C(SCPU_CTRL_SPI_CCT_IS_SHIFT), 
        .D(N363), .Y(N373) );
  CLKBUFX2TF U307 ( .A(\SCPU_CTRL_SPI_IO_CONTROL[6] ), .Y(N291) );
  NOR3X4TF U308 ( .A(N350), .B(N349), .C(N293), .Y(N361) );
  NAND2X1TF U309 ( .A(N424), .B(SCPU_CTRL_SPI_PUT_IS_ADDR_LEN_NZ), .Y(N414) );
  NOR2X1TF U310 ( .A(N336), .B(N352), .Y(N348) );
  NAND2X1TF U311 ( .A(I_CTRL_BGN), .B(N323), .Y(N331) );
  NOR2X1TF U312 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[3] ), .B(N296), .Y(N167)
         );
  AOI222XLTF U313 ( .A0(N361), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[1]), .B0(N360), 
        .B1(Q_FROM_SRAM[1]), .C0(N359), .C1(SCPU_CTRL_SPI_PUT_SRAM_REGS[2]), 
        .Y(N353) );
  AOI222XLTF U314 ( .A0(N361), .A1(I_SPI_SO), .B0(N360), .B1(Q_FROM_SRAM[0]), 
        .C0(SCPU_CTRL_SPI_PUT_SRAM_REGS[1]), .C1(N359), .Y(N362) );
  AOI222XLTF U315 ( .A0(N361), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[3]), .B0(N360), 
        .B1(Q_FROM_SRAM[3]), .C0(N359), .C1(SCPU_CTRL_SPI_PUT_SRAM_REGS[4]), 
        .Y(N355) );
  AOI222XLTF U316 ( .A0(N361), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[2]), .B0(N360), 
        .B1(Q_FROM_SRAM[2]), .C0(N359), .C1(SCPU_CTRL_SPI_PUT_SRAM_REGS[3]), 
        .Y(N354) );
  AOI222XLTF U317 ( .A0(N361), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[5]), .B0(N360), 
        .B1(Q_FROM_SRAM[5]), .C0(N359), .C1(SCPU_CTRL_SPI_PUT_SRAM_REGS[6]), 
        .Y(N357) );
  AOI222XLTF U318 ( .A0(N361), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[4]), .B0(N360), 
        .B1(Q_FROM_SRAM[4]), .C0(N359), .C1(SCPU_CTRL_SPI_PUT_SRAM_REGS[5]), 
        .Y(N356) );
  AOI222XLTF U319 ( .A0(N361), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[6]), .B0(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[7]), .B1(N359), .C0(N360), .C1(
        Q_FROM_SRAM[6]), .Y(N358) );
  NAND3X1TF U320 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .B(
        \SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .C(N103), .Y(N351) );
  NAND2X1TF U321 ( .A(N319), .B(N318), .Y(A_AFTER_MUX[8]) );
  NAND2X1TF U322 ( .A(N314), .B(N313), .Y(A_AFTER_MUX[7]) );
  NAND2X1TF U323 ( .A(N312), .B(N311), .Y(A_AFTER_MUX[6]) );
  NAND2X1TF U324 ( .A(N310), .B(N309), .Y(A_AFTER_MUX[5]) );
  NAND2X1TF U325 ( .A(N308), .B(N307), .Y(A_AFTER_MUX[4]) );
  NAND2X1TF U326 ( .A(N306), .B(N305), .Y(A_AFTER_MUX[3]) );
  NAND2X1TF U327 ( .A(N304), .B(N303), .Y(A_AFTER_MUX[2]) );
  NAND2X1TF U328 ( .A(N302), .B(N301), .Y(A_AFTER_MUX[1]) );
  CLKBUFX2TF U329 ( .A(N417), .Y(N292) );
  INVX2TF U330 ( .A(N291), .Y(N417) );
  AO21X1TF U331 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[3] ), .A1(N296), .B0(
        N167), .Y(SCPU_CTRL_SPI_CCT_N53) );
  NAND2X1TF U332 ( .A(N424), .B(N418), .Y(N420) );
  NOR2X1TF U333 ( .A(N350), .B(N348), .Y(N385) );
  NOR2X1TF U334 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ), .B(N297), .Y(N298)
         );
  NAND2X1TF U335 ( .A(N284), .B(N326), .Y(N297) );
  NOR2X1TF U336 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ), .B(N327), .Y(N326)
         );
  INVX2TF U337 ( .A(N331), .Y(N161) );
  NAND2X1TF U338 ( .A(N167), .B(N168), .Y(N323) );
  OR3X1TF U339 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ), .B(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ), .C(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .Y(N296) );
  NOR2X2TF U340 ( .A(N293), .B(N352), .Y(N359) );
  NAND3X1TF U341 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .B(N273), .C(N271), 
        .Y(N352) );
  OAI2BB2XLTF U342 ( .B0(N339), .B1(N414), .A0N(
        \SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .A1N(N335), .Y(N213) );
  OAI2BB1X1TF U343 ( .A0N(N320), .A1N(\SCPU_CTRL_SPI_CCT_REG_BITS[8] ), .B0(
        N299), .Y(A_AFTER_MUX[0]) );
  OAI221XLTF U344 ( .A0(N105), .A1(SCPU_CTRL_SPI_A_SPI[0]), .B0(N300), .B1(
        SCPU_CTRL_SPI_I_ADDR[0]), .C0(N264), .Y(N299) );
  AO22X1TF U345 ( .A0(N321), .A1(I_CTRL_SO), .B0(SCPU_CTRL_SPI_D_DATAOUT[0]), 
        .B1(N263), .Y(D_AFTER_MUX[0]) );
  NOR2X1TF U346 ( .A(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ), .B(N334), .Y(N336)
         );
  NAND2X1TF U347 ( .A(N268), .B(N279), .Y(N222) );
  NOR2X2TF U348 ( .A(N374), .B(N300), .Y(N317) );
  NOR2X2TF U349 ( .A(N300), .B(N382), .Y(N315) );
  NAND2X2TF U350 ( .A(SCPU_CTRL_SPI_IS_I_ADDR), .B(N263), .Y(N382) );
  NOR2X2TF U351 ( .A(I_CTRL_BGN), .B(N105), .Y(N316) );
  CLKBUFX2TF U352 ( .A(N292), .Y(N294) );
  AO21X1TF U353 ( .A0(\SCPU_CTRL_SPI_IO_DATAOUTA[6] ), .A1(N417), .B0(N396), 
        .Y(N87) );
  AO22X1TF U354 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[4]), .B0(N384), .B1(I_ADC_PI[4]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[4]) );
  AO22X1TF U355 ( .A0(N265), .A1(SCPU_CTRL_SPI_FOUT[8]), .B0(N384), .B1(
        I_ADC_PI[8]), .Y(SCPU_CTRL_SPI_IO_DATAINA[8]) );
  AO22X1TF U356 ( .A0(N265), .A1(SCPU_CTRL_SPI_FOUT[9]), .B0(N384), .B1(
        I_ADC_PI[9]), .Y(SCPU_CTRL_SPI_IO_DATAINA[9]) );
  AO22X1TF U357 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[7]), .B0(N384), .B1(I_ADC_PI[7]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[7]) );
  AO22X1TF U358 ( .A0(N265), .A1(SCPU_CTRL_SPI_FOUT[6]), .B0(N384), .B1(
        I_ADC_PI[6]), .Y(SCPU_CTRL_SPI_IO_DATAINA[6]) );
  INVX2TF U359 ( .A(N265), .Y(N384) );
  AOI31X1TF U360 ( .A0(N424), .A1(N423), .A2(N274), .B0(N280), .Y(N46) );
  NOR2X1TF U361 ( .A(\SCPU_CTRL_SPI_PUT_CNT_STATE[0] ), .B(N388), .Y(
        SCPU_CTRL_SPI_PUT_N108) );
  OAI32X1TF U362 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ), .A1(
        \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .A2(N420), .B0(N421), .B1(N277), 
        .Y(N37) );
  AOI32X1TF U363 ( .A0(N424), .A1(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] ), .A2(
        N423), .B0(N422), .B1(N274), .Y(N43) );
  AOI32X1TF U364 ( .A0(N421), .A1(N422), .A2(N277), .B0(N286), .B1(N422), .Y(
        N40) );
  OAI211X1TF U365 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] ), .A1(
        \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[4] ), .B0(N424), .C0(N423), .Y(N422)
         );
  NOR2X1TF U366 ( .A(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .B(N419), .Y(N421)
         );
  OAI211X1TF U367 ( .A0(N348), .A1(N278), .B0(N351), .C0(N347), .Y(N208) );
  OAI211X1TF U368 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .A1(N347), .B0(
        N351), .C0(N346), .Y(N209) );
  OAI21X1TF U369 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .A1(N385), .B0(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .Y(N346) );
  OAI31X1TF U370 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .A1(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .A2(N385), .B0(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ), .Y(N345) );
  AOI22X1TF U371 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ), .A1(N343), .B0(
        N344), .B1(N287), .Y(N211) );
  AOI21X1TF U372 ( .A0(N349), .A1(N334), .B0(N385), .Y(N343) );
  INVX2TF U373 ( .A(N385), .Y(N387) );
  OAI21X1TF U374 ( .A0(N326), .A1(N284), .B0(N297), .Y(SCPU_CTRL_SPI_CCT_N55)
         );
  OAI22X1TF U375 ( .A0(I_CTRL_MODE[0]), .A1(N329), .B0(N328), .B1(N331), .Y(
        N218) );
  AOI21X1TF U376 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ), .A1(N327), .B0(
        N326), .Y(N328) );
  INVX2TF U377 ( .A(N167), .Y(N327) );
  OAI21X1TF U378 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .A1(N331), .B0(
        N330), .Y(N217) );
  NOR4X1TF U379 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[7] ), .B(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ), .C(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[5] ), .D(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ), .Y(N168) );
  INVX2TF U380 ( .A(N353), .Y(N206) );
  INVX2TF U381 ( .A(N362), .Y(N200) );
  INVX2TF U382 ( .A(N355), .Y(N204) );
  INVX2TF U383 ( .A(N354), .Y(N205) );
  INVX2TF U384 ( .A(N357), .Y(N202) );
  INVX2TF U385 ( .A(N356), .Y(N203) );
  INVX2TF U386 ( .A(N358), .Y(N201) );
  INVX2TF U387 ( .A(N352), .Y(N349) );
  INVX2TF U388 ( .A(N351), .Y(N350) );
  OAI21X1TF U389 ( .A0(N376), .A1(N373), .B0(N365), .Y(N198) );
  AOI22X1TF U390 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[2] ), .A1(N266), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[1] ), .B1(N371), .Y(N365) );
  OAI21X1TF U391 ( .A0(N377), .A1(N373), .B0(N366), .Y(N197) );
  AOI22X1TF U392 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[3] ), .A1(N266), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[2] ), .B1(N371), .Y(N366) );
  OAI21X1TF U393 ( .A0(N381), .A1(N373), .B0(N370), .Y(N193) );
  AOI22X1TF U394 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[7] ), .A1(N266), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[6] ), .B1(N371), .Y(N370) );
  OAI21X1TF U395 ( .A0(N380), .A1(N373), .B0(N369), .Y(N194) );
  AOI22X1TF U396 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[6] ), .A1(N266), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[5] ), .B1(N371), .Y(N369) );
  OAI21X1TF U397 ( .A0(N378), .A1(N373), .B0(N367), .Y(N196) );
  AOI22X1TF U398 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[4] ), .A1(N266), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[3] ), .B1(N371), .Y(N367) );
  OAI21X1TF U399 ( .A0(N383), .A1(N373), .B0(N372), .Y(N192) );
  AOI22X1TF U400 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[8] ), .A1(N266), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[7] ), .B1(N371), .Y(N372) );
  OAI21X1TF U401 ( .A0(N379), .A1(N373), .B0(N368), .Y(N195) );
  AOI22X1TF U402 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[5] ), .A1(N266), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[4] ), .B1(N371), .Y(N368) );
  OAI21X1TF U403 ( .A0(N375), .A1(N373), .B0(N364), .Y(N199) );
  AOI22X1TF U404 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[1] ), .A1(N266), .B0(
        I_CTRL_SO), .B1(N371), .Y(N364) );
  OAI211X4TF U405 ( .A0(N95), .A1(N363), .B0(N268), .C0(
        SCPU_CTRL_SPI_CCT_IS_SHIFT), .Y(N371) );
  INVX2TF U406 ( .A(I_CTRL_MODE[1]), .Y(N363) );
  AND2X2TF U407 ( .A(N338), .B(N271), .Y(N225) );
  NOR2X1TF U408 ( .A(N95), .B(N268), .Y(N223) );
  AND2X2TF U409 ( .A(SCPU_CTRL_SPI_CEN), .B(I_CTRL_BGN), .Y(CEN_AFTER_MUX) );
  AOI32X1TF U410 ( .A0(N105), .A1(N264), .A2(SCPU_CTRL_SPI_D_WE), .B0(
        I_CTRL_BGN), .B1(N281), .Y(WEN_AFTER_MUX) );
  NOR2X1TF U411 ( .A(N379), .B(N382), .Y(SCPU_CTRL_SPI_I_DATAIN[4]) );
  NOR2X1TF U412 ( .A(N375), .B(N382), .Y(SCPU_CTRL_SPI_I_DATAIN[0]) );
  NOR2X1TF U413 ( .A(N376), .B(N382), .Y(SCPU_CTRL_SPI_I_DATAIN[1]) );
  NOR2X1TF U414 ( .A(N380), .B(N382), .Y(SCPU_CTRL_SPI_I_DATAIN[5]) );
  NOR2X1TF U415 ( .A(N377), .B(N382), .Y(SCPU_CTRL_SPI_I_DATAIN[2]) );
  NOR2X1TF U416 ( .A(N381), .B(N382), .Y(SCPU_CTRL_SPI_I_DATAIN[6]) );
  NOR2X1TF U417 ( .A(N378), .B(N382), .Y(SCPU_CTRL_SPI_I_DATAIN[3]) );
  NOR2X1TF U418 ( .A(N383), .B(N382), .Y(SCPU_CTRL_SPI_I_DATAIN[7]) );
  NOR2X1TF U419 ( .A(N378), .B(N374), .Y(SCPU_CTRL_SPI_D_DATAIN[3]) );
  INVX2TF U420 ( .A(Q_FROM_SRAM[3]), .Y(N378) );
  NOR2X1TF U421 ( .A(N377), .B(N374), .Y(SCPU_CTRL_SPI_D_DATAIN[2]) );
  INVX2TF U422 ( .A(Q_FROM_SRAM[2]), .Y(N377) );
  NOR2X1TF U423 ( .A(N381), .B(N374), .Y(SCPU_CTRL_SPI_D_DATAIN[6]) );
  INVX2TF U424 ( .A(Q_FROM_SRAM[6]), .Y(N381) );
  NOR2X1TF U425 ( .A(N379), .B(N374), .Y(SCPU_CTRL_SPI_D_DATAIN[4]) );
  INVX2TF U426 ( .A(Q_FROM_SRAM[4]), .Y(N379) );
  NOR2X1TF U427 ( .A(N375), .B(N374), .Y(SCPU_CTRL_SPI_D_DATAIN[0]) );
  INVX2TF U428 ( .A(Q_FROM_SRAM[0]), .Y(N375) );
  NOR2X1TF U429 ( .A(N376), .B(N374), .Y(SCPU_CTRL_SPI_D_DATAIN[1]) );
  INVX2TF U430 ( .A(Q_FROM_SRAM[1]), .Y(N376) );
  NOR2X1TF U431 ( .A(N383), .B(N374), .Y(SCPU_CTRL_SPI_D_DATAIN[7]) );
  INVX2TF U432 ( .A(Q_FROM_SRAM[7]), .Y(N383) );
  NOR2X1TF U433 ( .A(N380), .B(N374), .Y(SCPU_CTRL_SPI_D_DATAIN[5]) );
  INVX2TF U434 ( .A(Q_FROM_SRAM[5]), .Y(N380) );
  OAI32X1TF U435 ( .A0(N293), .A1(N105), .A2(N332), .B0(N419), .B1(N293), .Y(
        N216) );
  INVX2TF U436 ( .A(N424), .Y(N419) );
  OAI21X1TF U437 ( .A0(N103), .A1(N341), .B0(N340), .Y(N212) );
  OAI32X1TF U438 ( .A0(N339), .A1(N411), .A2(N338), .B0(
        \SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .B1(N337), .Y(N340) );
  NOR2X1TF U439 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .B(
        \SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .Y(N338) );
  AOI21X1TF U440 ( .A0(N336), .A1(N337), .B0(\SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), 
        .Y(N341) );
  INVX2TF U441 ( .A(N339), .Y(N337) );
  AOI21X1TF U442 ( .A0(N271), .A1(N333), .B0(N388), .Y(N339) );
  NOR3X1TF U443 ( .A(\SCPU_CTRL_SPI_PUT_CNT_STATE[0] ), .B(
        \SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .C(\SCPU_CTRL_SPI_PUT_CNT_STATE[2] ), .Y(N388) );
  INVX2TF U444 ( .A(N342), .Y(N334) );
  NOR3X1TF U445 ( .A(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ), .B(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .C(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .Y(N342) );
  AOI22X1TF U446 ( .A0(SCPU_CTRL_SPI_A_SPI[8]), .A1(N316), .B0(N315), .B1(
        SCPU_CTRL_SPI_I_ADDR[8]), .Y(N319) );
  AOI22X1TF U447 ( .A0(SCPU_CTRL_SPI_A_SPI[7]), .A1(N316), .B0(N315), .B1(
        SCPU_CTRL_SPI_I_ADDR[7]), .Y(N314) );
  AOI22X1TF U448 ( .A0(SCPU_CTRL_SPI_A_SPI[6]), .A1(N316), .B0(N315), .B1(
        SCPU_CTRL_SPI_I_ADDR[6]), .Y(N312) );
  AOI22X1TF U449 ( .A0(SCPU_CTRL_SPI_A_SPI[5]), .A1(N316), .B0(N315), .B1(
        SCPU_CTRL_SPI_I_ADDR[5]), .Y(N310) );
  AOI22X1TF U450 ( .A0(SCPU_CTRL_SPI_A_SPI[4]), .A1(N316), .B0(N315), .B1(
        SCPU_CTRL_SPI_I_ADDR[4]), .Y(N308) );
  AOI22X1TF U451 ( .A0(SCPU_CTRL_SPI_A_SPI[3]), .A1(N316), .B0(N315), .B1(
        SCPU_CTRL_SPI_I_ADDR[3]), .Y(N306) );
  AOI22X1TF U452 ( .A0(SCPU_CTRL_SPI_A_SPI[2]), .A1(N316), .B0(N315), .B1(
        SCPU_CTRL_SPI_I_ADDR[2]), .Y(N304) );
  AOI22X1TF U453 ( .A0(SCPU_CTRL_SPI_A_SPI[1]), .A1(N316), .B0(N315), .B1(
        SCPU_CTRL_SPI_I_ADDR[1]), .Y(N302) );
  OAI31X1TF U454 ( .A0(SCPU_CTRL_SPI_A_SPI[2]), .A1(N416), .A2(N410), .B0(N409), .Y(N83) );
  AOI22X1TF U455 ( .A0(SCPU_CTRL_SPI_A_SPI[2]), .A1(N408), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[2] ), .B1(N293), .Y(N409) );
  AOI31X1TF U456 ( .A0(N411), .A1(SCPU_CTRL_SPI_A_SPI[0]), .A2(
        SCPU_CTRL_SPI_A_SPI[1]), .B0(N294), .Y(N408) );
  OAI31X1TF U457 ( .A0(SCPU_CTRL_SPI_A_SPI[1]), .A1(N416), .A2(N285), .B0(N413), .Y(N82) );
  AOI22X1TF U458 ( .A0(SCPU_CTRL_SPI_A_SPI[1]), .A1(N412), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[1] ), .B1(N293), .Y(N413) );
  AOI21X1TF U459 ( .A0(N411), .A1(SCPU_CTRL_SPI_A_SPI[0]), .B0(N294), .Y(N412)
         );
  OAI31X1TF U460 ( .A0(SCPU_CTRL_SPI_A_SPI[3]), .A1(N416), .A2(N407), .B0(N406), .Y(N84) );
  AOI22X1TF U461 ( .A0(SCPU_CTRL_SPI_A_SPI[3]), .A1(N405), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[3] ), .B1(N294), .Y(N406) );
  AOI21X1TF U462 ( .A0(N411), .A1(N404), .B0(N294), .Y(N405) );
  OAI31X1TF U463 ( .A0(SCPU_CTRL_SPI_A_SPI[4]), .A1(N416), .A2(N403), .B0(N402), .Y(N85) );
  AOI22X1TF U464 ( .A0(SCPU_CTRL_SPI_A_SPI[4]), .A1(N401), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[4] ), .B1(N294), .Y(N402) );
  AOI31X1TF U465 ( .A0(N411), .A1(N404), .A2(SCPU_CTRL_SPI_A_SPI[3]), .B0(N294), .Y(N401) );
  OAI21X1TF U466 ( .A0(SCPU_CTRL_SPI_A_SPI[0]), .A1(N416), .B0(N415), .Y(N81)
         );
  AOI32X1TF U467 ( .A0(SCPU_CTRL_SPI_A_SPI[0]), .A1(N291), .A2(N414), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[0] ), .B1(N293), .Y(N415) );
  OAI21X1TF U468 ( .A0(SCPU_CTRL_SPI_A_SPI[5]), .A1(N400), .B0(N399), .Y(N86)
         );
  AOI22X1TF U469 ( .A0(SCPU_CTRL_SPI_A_SPI[5]), .A1(N398), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[5] ), .B1(N294), .Y(N399) );
  OAI31X1TF U470 ( .A0(SCPU_CTRL_SPI_A_SPI[8]), .A1(N283), .A2(N392), .B0(N391), .Y(N89) );
  AOI22X1TF U471 ( .A0(SCPU_CTRL_SPI_A_SPI[8]), .A1(N390), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[8] ), .B1(N293), .Y(N391) );
  OAI21X1TF U472 ( .A0(SCPU_CTRL_SPI_A_SPI[7]), .A1(N416), .B0(N394), .Y(N390)
         );
  OAI21X1TF U473 ( .A0(N394), .A1(N283), .B0(N393), .Y(N88) );
  NOR3X1TF U474 ( .A(N397), .B(N276), .C(N282), .Y(N389) );
  OAI32X1TF U475 ( .A0(SCPU_CTRL_SPI_A_SPI[6]), .A1(N276), .A2(N400), .B0(N395), .B1(N282), .Y(N396) );
  OAI31X1TF U476 ( .A0(N414), .A1(N397), .A2(N276), .B0(N291), .Y(N395) );
  OR2X2TF U477 ( .A(N397), .B(N416), .Y(N400) );
  NAND2X2TF U478 ( .A(N291), .B(N411), .Y(N416) );
  INVX2TF U479 ( .A(N414), .Y(N411) );
  AND3X2TF U480 ( .A(N289), .B(\SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .C(N103), 
        .Y(N424) );
  INVX2TF U481 ( .A(N407), .Y(N404) );
  AND2X2TF U482 ( .A(N332), .B(N271), .Y(N224) );
  NOR2X1TF U483 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .B(N273), .Y(N332) );
  NOR3X1TF U484 ( .A(N105), .B(N275), .C(N272), .Y(I_SCLK1) );
  NOR3X1TF U485 ( .A(\SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .B(N105), .C(N272), 
        .Y(I_SCLK2) );
  OAI2BB1X1TF U486 ( .A0N(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .A1N(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ), .B0(N295), .Y(
        SCPU_CTRL_SPI_CCT_N51) );
  OAI2BB1X1TF U487 ( .A0N(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ), .A1N(N295), 
        .B0(N296), .Y(SCPU_CTRL_SPI_CCT_N52) );
  AO21X1TF U488 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ), .A1(N297), .B0(
        N298), .Y(SCPU_CTRL_SPI_CCT_N56) );
  XOR2X1TF U489 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[7] ), .B(N298), .Y(
        SCPU_CTRL_SPI_CCT_N57) );
  AO22X1TF U490 ( .A0(N321), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[1] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[1]), .B1(N264), .Y(D_AFTER_MUX[1]) );
  AO22X1TF U491 ( .A0(N321), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[2] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[2]), .B1(N264), .Y(D_AFTER_MUX[2]) );
  AO22X1TF U492 ( .A0(N321), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[3] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[3]), .B1(N264), .Y(D_AFTER_MUX[3]) );
  AO22X1TF U493 ( .A0(N321), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[4] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[4]), .B1(N264), .Y(D_AFTER_MUX[4]) );
  AO22X1TF U494 ( .A0(N321), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[5] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[5]), .B1(N264), .Y(D_AFTER_MUX[5]) );
  AO22X1TF U495 ( .A0(N321), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[6] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[6]), .B1(N264), .Y(D_AFTER_MUX[6]) );
  AO22X1TF U496 ( .A0(N321), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[7] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[7]), .B1(N264), .Y(D_AFTER_MUX[7]) );
  NAND2BX1TF U497 ( .AN(N222), .B(I_CTRL_MODE[1]), .Y(N221) );
  OAI221XLTF U498 ( .A0(N268), .A1(I_LOAD_N), .B0(N288), .B1(N323), .C0(
        I_CTRL_BGN), .Y(N322) );
  AO22X1TF U499 ( .A0(N268), .A1(N161), .B0(N325), .B1(N322), .Y(N219) );
  NAND3BX1TF U500 ( .AN(I_LOAD_N), .B(N325), .C(N324), .Y(N329) );
  AO21X1TF U501 ( .A0(I_CTRL_MODE[0]), .A1(I_CTRL_MODE[1]), .B0(N329), .Y(N330) );
  NAND2X1TF U502 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .B(N273), .Y(N333) );
  NAND2X1TF U503 ( .A(N342), .B(N348), .Y(N344) );
  NAND3X1TF U504 ( .A(N351), .B(N345), .C(N344), .Y(N210) );
  NAND2X1TF U505 ( .A(N348), .B(N278), .Y(N347) );
  AO22X1TF U506 ( .A0(N361), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[7]), .B0(
        Q_FROM_SRAM[7]), .B1(N360), .Y(N207) );
  AO22X1TF U507 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[0]), .B0(N384), .B1(I_ADC_PI[0]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[0]) );
  AO22X1TF U508 ( .A0(N265), .A1(SCPU_CTRL_SPI_FOUT[1]), .B0(N384), .B1(
        I_ADC_PI[1]), .Y(SCPU_CTRL_SPI_IO_DATAINA[1]) );
  AO22X1TF U509 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[2]), .B0(N384), .B1(I_ADC_PI[2]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[2]) );
  AO22X1TF U510 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[3]), .B0(N384), .B1(I_ADC_PI[3]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[3]) );
  AO22X1TF U511 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[5]), .B0(N384), .B1(I_ADC_PI[5]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[5]) );
  AO22X1TF U512 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .A1(
        \SCPU_CTRL_SPI_PUT_CNT_STATE[0] ), .B0(N275), .B1(
        SCPU_CTRL_SPI_PUT_N108), .Y(SCPU_CTRL_SPI_PUT_N109) );
  AO22X1TF U513 ( .A0(N388), .A1(N387), .B0(\SCPU_CTRL_SPI_PUT_CNT_STATE[2] ), 
        .B1(N386), .Y(SCPU_CTRL_SPI_PUT_N110) );
  NAND3X1TF U514 ( .A(N280), .B(N274), .C(N423), .Y(N418) );
  NAND3X1TF U515 ( .A(SCPU_CTRL_SPI_A_SPI[2]), .B(SCPU_CTRL_SPI_A_SPI[0]), .C(
        SCPU_CTRL_SPI_A_SPI[1]), .Y(N407) );
  NAND3X1TF U516 ( .A(SCPU_CTRL_SPI_A_SPI[4]), .B(N404), .C(
        SCPU_CTRL_SPI_A_SPI[3]), .Y(N397) );
  NAND2BX1TF U517 ( .AN(N416), .B(N389), .Y(N392) );
  AO21X1TF U518 ( .A0(N411), .A1(N389), .B0(N417), .Y(N394) );
  AOI2BB2X1TF U519 ( .B0(\SCPU_CTRL_SPI_IO_DATAOUTA[7] ), .B1(N293), .A0N(
        SCPU_CTRL_SPI_A_SPI[7]), .A1N(N392), .Y(N393) );
  AOI2BB1X1TF U520 ( .A0N(N414), .A1N(N397), .B0(N292), .Y(N398) );
  XNOR2X1TF U522 ( .A(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .B(N420), .Y(N34)
         );
endmodule

