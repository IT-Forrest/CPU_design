
module SHARE_SUPERALU_VG ( CLK, RST_N, X_IN, Y_IN, ALU_START, ALU_TYPE, MODE_TYPE, 
        OFFSET, FOUT, POUT, ALU_IS_DONE );
  input [12:0] X_IN;
  input [12:0] Y_IN;
  input [2:0] ALU_TYPE;
  input [1:0] MODE_TYPE;
  input [9:0] OFFSET;
  output [12:0] FOUT;
  output [12:0] POUT;
  input CLK, RST_N, ALU_START;
  output ALU_IS_DONE;
  wire   POST_WORK, PRE_WORK, \INDEX[2] , \RSHT_BITS[3] , SIGN_Y, C152_DATA4_0,
         C152_DATA4_1, C152_DATA4_2, C152_DATA4_3, C152_DATA4_4, C152_DATA4_5,
         C152_DATA4_6, C152_DATA4_7, C152_DATA4_8, C152_DATA4_9, C152_DATA4_10,
         C152_DATA4_11, N73, N74, N90, N91, N92, N121, N122, N123, N124, N128,
         N129, N657, N658, N659, N660, N661, N662, N663, N664, N665, N666,
         N667, N668, N669, N670, N671, N672, N673, N674, N675, N676, N677,
         N678, N679, N680, N681, N682, N683, N684, N685, N686, N687, N688,
         N689, N690, N691, N692, N693, N694, N695, N696, N697, N698, N699,
         N700, N701, N702, N703, N704, N705, N706, N707, N708, N709, N710,
         N711, N712, N713, N714, N715, N716, N717, N718, N719, N720, N721,
         N722, N723, N724, N725, N726, C2_Z_11, C2_Z_10, C2_Z_9, C2_Z_8,
         C2_Z_7, C2_Z_6, C2_Z_5, C2_Z_4, C2_Z_3, C2_Z_2, C2_Z_1, C2_Z_0,
         DP_OP_333_124_4748_N57, DP_OP_333_124_4748_N29,
         DP_OP_333_124_4748_N28, DP_OP_333_124_4748_N27,
         DP_OP_333_124_4748_N26, DP_OP_333_124_4748_N25,
         DP_OP_333_124_4748_N24, DP_OP_333_124_4748_N23,
         DP_OP_333_124_4748_N22, DP_OP_333_124_4748_N21,
         DP_OP_333_124_4748_N20, DP_OP_333_124_4748_N19,
         DP_OP_333_124_4748_N18, DP_OP_333_124_4748_N12,
         DP_OP_333_124_4748_N11, DP_OP_333_124_4748_N10, DP_OP_333_124_4748_N9,
         DP_OP_333_124_4748_N8, DP_OP_333_124_4748_N7, DP_OP_333_124_4748_N6,
         DP_OP_333_124_4748_N5, DP_OP_333_124_4748_N4, DP_OP_333_124_4748_N3,
         DP_OP_333_124_4748_N2, DP_OP_333_124_4748_N1, INTADD_0_CI,
         \INTADD_0_SUM[6] , \INTADD_0_SUM[5] , \INTADD_0_SUM[4] ,
         \INTADD_0_SUM[3] , \INTADD_0_SUM[2] , \INTADD_0_SUM[1] ,
         \INTADD_0_SUM[0] , INTADD_0_N7, INTADD_0_N6, INTADD_0_N5, INTADD_0_N4,
         INTADD_0_N3, INTADD_0_N2, INTADD_0_N1, ADD_X_132_1_N13,
         ADD_X_132_1_N12, ADD_X_132_1_N11, ADD_X_132_1_N10, ADD_X_132_1_N9,
         ADD_X_132_1_N8, ADD_X_132_1_N7, ADD_X_132_1_N6, ADD_X_132_1_N5,
         ADD_X_132_1_N4, ADD_X_132_1_N3, ADD_X_132_1_N2, N1, N2, N3, N4, N5,
         N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N81,
         N82, N83, N84, N85, N86, N87, N88, N89, N93, N94, N95, N96, N97, N98,
         N99, N100, N101, N102, N103, N104, N105, N106, N107, N108, N109, N110,
         N111, N112, N113, N114, N115, N116, N117, N118, N119, N120, N125,
         N126, N127, N130, N131, N132, N133, N134, N135, N136, N137, N138,
         N139, N140, N141, N142, N143, N144, N145, N146, N147, N149, N150,
         N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161,
         N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172,
         N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183,
         N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194,
         N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205,
         N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216,
         N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227,
         N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238,
         N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249,
         N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260,
         N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271,
         N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282,
         N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293,
         N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304,
         N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315,
         N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326,
         N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337,
         N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, N348,
         N349, N350, N351, N352, N353, N354, N355, N356, N357, N358, N359,
         N360, N361, N362, N363, N364, N365, N366, N367, N368, N369, N370,
         N371, N372, N373, N374, N375, N376, N377, N378, N379, N380, N381,
         N382, N383, N384, N385, N386, N387, N388, N389, N390, N391, N392,
         N393, N394, N395, N396, N397, N398, N399, N400, N401, N402, N403,
         N404, N405, N406, N407, N408, N409, N410, N411, N412, N413, N414,
         N415, N416, N417, N418, N419, N420, N421, N422, N423, N424, N425,
         N426, N427, N428, N429, N430, N431, N432, N433, N434, N435, N436,
         N437, N438, N439, N440, N441, N442, N443, N444, N445, N446, N447,
         N448, N449, N450, N451, N452, N453, N454, N455, N456, N457, N458,
         N459, N460, N461, N462, N463, N464, N465, N466, N467, N468, N469,
         N470, N471, N472, N473, N474, N475, N476, N477, N478, N479, N480,
         N481, N482, N483, N484, N485, N486, N487, N488, N489, N490, N491,
         N492, N493, N494, N495, N496, N497, N498, N499, N500, N501, N502,
         N503, N504, N505, N506, N507, N508, N509, N510, N511, N512, N513,
         N514, N515, N516, N517, N518, N519, N520, N521, N522, N523, N524,
         N525, N526, N527, N528, N529, N530, N531, N532, N533, N534, N535,
         N536, N537, N538, N539, N540, N541, N542, N543, N544, N545, N546,
         N547, N548, N549, N550, N551, N552, N553, N554, N555, N556, N557,
         N558, N559, N560, N561, N562, N563, N564, N565, N566, N567, N568,
         N569, N570, N571, N572, N573, N574, N575, N576, N577, N578, N579,
         N580, N581, N582, N583, N584, N585, N586, N587, N588, N589, N590,
         N591, N592, N593, N594, N595, N596, N597, N598, N599, N600, N601,
         N602, N603, N604, N605, N606, N607, N608, N609, N610, N611, N612,
         N613, N614, N615, N616, N617, N618, N619, N620, N621, N622, N623,
         N624, N625, N626, N627, N628, N629, N630, N631, N632, N633, N634,
         N635, N636, N637, N638, N639, N640, N641, N642, N643, N644, N645,
         N646, N647, N648, N649, N650, N651, N652, N653, N654, N655, N656,
         N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737,
         N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748,
         N749, N750, N751, N752, N753, N754, N755, N756, N757, N758, N759,
         N760, N761, N762, N763, N764, N765, N766, N767, N768, N769, N770,
         N771, N772, N773, N774, N775, N776, N777, N778, N779, N780, N781,
         N782, N783, N784, N785, N786, N787, N788, N789, N790, N791, N792,
         N793, N794, N795, N796, N797, N798, N799, N800, N801, N802, N803,
         N804, N805, N806, N807, N808, N809, N810, N811, N812, N813, N814,
         N815, N816, N817, N818, N819, N820, N821, N822, N823, N824, N825,
         N826, N827, N828, N829, N830, N831, N832, N833, N834, N835, N836,
         N837, N838, N839, N840, N841, N842, N843, N844, N845, N846, N847,
         N848, N849, N850, N851, N852, N853, N854, N855, N856, N857, N858,
         N859, N860, N861, N862, N863, N864, N865, N866, N867, N868, N869,
         N870, N871, N872, N873, N874, N875, N876, N877, N878, N879, N880,
         N881, N882, N883, N884, N885, N886, N887, N888, N889, N890, N891,
         N892, N893, N894, N895, N896, N897, N898, N899, N900, N901, N902,
         N903, N904, N905, N906, N907, N908, N909, N910, N911, N912, N913,
         N914, N915, N916, N917, N918, N919, N920, N921, N922, N923, N924,
         N925, N926, N927, N928, N929, N930, N931, N932, N933, N934, N935,
         N936, N937, N938, N939, N940, N941, N942, N943, N944, N945, N946,
         N947, N948, N949, N950, N951, N952, N953, N954, N955, N956, N957,
         N958, N959, N960, N961, N962, N963, N964, N965, N966, N967, N968,
         N969, N970, N971, N972, N973, N974, N975, N976, N977, N978, N979,
         N980, N981, N982, N983, N984, N985, N986, N987, N988, N989, N990,
         N991, N992, N993, N994, N995, N996, N997, N998, N999, N1000, N1001,
         N1002, N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011,
         N1012, N1013, N1014, N1015, N1016, N1017, N1018, N1019;
  wire   [12:9] XTEMP;
  wire   [12:0] DIVISION_HEAD;
  wire   [8:0] DIVISION_REMA;
  wire   [12:0] OPER_A;
  wire   [12:0] OPER_B;
  wire   [12:0] SUM_AB;
  wire   [12:0] ZTEMP;
  wire   [3:2] STEP;

  XOR2X1TF \DP_OP_333_124_4748/U28  ( .A(N81), .B(C2_Z_0), .Y(
        DP_OP_333_124_4748_N29) );
  XOR2X1TF \DP_OP_333_124_4748/U27  ( .A(N81), .B(C2_Z_1), .Y(
        DP_OP_333_124_4748_N28) );
  XOR2X1TF \DP_OP_333_124_4748/U26  ( .A(N81), .B(C2_Z_2), .Y(
        DP_OP_333_124_4748_N27) );
  XOR2X1TF \DP_OP_333_124_4748/U25  ( .A(N971), .B(C2_Z_3), .Y(
        DP_OP_333_124_4748_N26) );
  XOR2X1TF \DP_OP_333_124_4748/U24  ( .A(N81), .B(C2_Z_4), .Y(
        DP_OP_333_124_4748_N25) );
  XOR2X1TF \DP_OP_333_124_4748/U23  ( .A(N81), .B(C2_Z_5), .Y(
        DP_OP_333_124_4748_N24) );
  XOR2X1TF \DP_OP_333_124_4748/U22  ( .A(N81), .B(C2_Z_6), .Y(
        DP_OP_333_124_4748_N23) );
  XOR2X1TF \DP_OP_333_124_4748/U21  ( .A(N971), .B(C2_Z_7), .Y(
        DP_OP_333_124_4748_N22) );
  XOR2X1TF \DP_OP_333_124_4748/U20  ( .A(N81), .B(C2_Z_8), .Y(
        DP_OP_333_124_4748_N21) );
  XOR2X1TF \DP_OP_333_124_4748/U19  ( .A(N971), .B(C2_Z_9), .Y(
        DP_OP_333_124_4748_N20) );
  XOR2X1TF \DP_OP_333_124_4748/U18  ( .A(N81), .B(C2_Z_10), .Y(
        DP_OP_333_124_4748_N19) );
  XOR2X1TF \DP_OP_333_124_4748/U17  ( .A(N971), .B(C2_Z_11), .Y(
        DP_OP_333_124_4748_N18) );
  CMPR32X2TF \DP_OP_333_124_4748/U13  ( .A(DP_OP_333_124_4748_N57), .B(N971), 
        .C(DP_OP_333_124_4748_N29), .CO(DP_OP_333_124_4748_N12), .S(
        C152_DATA4_0) );
  ADDHXLTF \DP_OP_333_124_4748/U12  ( .A(DP_OP_333_124_4748_N28), .B(
        DP_OP_333_124_4748_N12), .CO(DP_OP_333_124_4748_N11), .S(C152_DATA4_1)
         );
  ADDHXLTF \DP_OP_333_124_4748/U11  ( .A(DP_OP_333_124_4748_N27), .B(
        DP_OP_333_124_4748_N11), .CO(DP_OP_333_124_4748_N10), .S(C152_DATA4_2)
         );
  ADDHXLTF \DP_OP_333_124_4748/U10  ( .A(DP_OP_333_124_4748_N26), .B(
        DP_OP_333_124_4748_N10), .CO(DP_OP_333_124_4748_N9), .S(C152_DATA4_3)
         );
  ADDHXLTF \DP_OP_333_124_4748/U9  ( .A(DP_OP_333_124_4748_N25), .B(
        DP_OP_333_124_4748_N9), .CO(DP_OP_333_124_4748_N8), .S(C152_DATA4_4)
         );
  ADDHXLTF \DP_OP_333_124_4748/U8  ( .A(DP_OP_333_124_4748_N24), .B(
        DP_OP_333_124_4748_N8), .CO(DP_OP_333_124_4748_N7), .S(C152_DATA4_5)
         );
  ADDHXLTF \DP_OP_333_124_4748/U7  ( .A(DP_OP_333_124_4748_N23), .B(
        DP_OP_333_124_4748_N7), .CO(DP_OP_333_124_4748_N6), .S(C152_DATA4_6)
         );
  ADDHXLTF \DP_OP_333_124_4748/U6  ( .A(DP_OP_333_124_4748_N22), .B(
        DP_OP_333_124_4748_N6), .CO(DP_OP_333_124_4748_N5), .S(C152_DATA4_7)
         );
  ADDHXLTF \DP_OP_333_124_4748/U5  ( .A(DP_OP_333_124_4748_N21), .B(
        DP_OP_333_124_4748_N5), .CO(DP_OP_333_124_4748_N4), .S(C152_DATA4_8)
         );
  ADDHXLTF \DP_OP_333_124_4748/U4  ( .A(DP_OP_333_124_4748_N20), .B(
        DP_OP_333_124_4748_N4), .CO(DP_OP_333_124_4748_N3), .S(C152_DATA4_9)
         );
  ADDHXLTF \DP_OP_333_124_4748/U3  ( .A(DP_OP_333_124_4748_N19), .B(
        DP_OP_333_124_4748_N3), .CO(DP_OP_333_124_4748_N2), .S(C152_DATA4_10)
         );
  ADDHXLTF \DP_OP_333_124_4748/U2  ( .A(DP_OP_333_124_4748_N18), .B(
        DP_OP_333_124_4748_N2), .CO(DP_OP_333_124_4748_N1), .S(C152_DATA4_11)
         );
  CMPR32X2TF \intadd_0/U8  ( .A(X_IN[1]), .B(DIVISION_HEAD[5]), .C(INTADD_0_CI), .CO(INTADD_0_N7), .S(\INTADD_0_SUM[0] ) );
  CMPR32X2TF \intadd_0/U7  ( .A(X_IN[2]), .B(DIVISION_HEAD[6]), .C(INTADD_0_N7), .CO(INTADD_0_N6), .S(\INTADD_0_SUM[1] ) );
  CMPR32X2TF \intadd_0/U6  ( .A(N94), .B(DIVISION_HEAD[7]), .C(INTADD_0_N6), 
        .CO(INTADD_0_N5), .S(\INTADD_0_SUM[2] ) );
  CMPR32X2TF \intadd_0/U5  ( .A(X_IN[4]), .B(DIVISION_HEAD[8]), .C(INTADD_0_N5), .CO(INTADD_0_N4), .S(\INTADD_0_SUM[3] ) );
  CMPR32X2TF \intadd_0/U4  ( .A(N106), .B(DIVISION_HEAD[9]), .C(INTADD_0_N4), 
        .CO(INTADD_0_N3), .S(\INTADD_0_SUM[4] ) );
  CMPR32X2TF \intadd_0/U3  ( .A(X_IN[6]), .B(DIVISION_HEAD[10]), .C(
        INTADD_0_N3), .CO(INTADD_0_N2), .S(\INTADD_0_SUM[5] ) );
  CMPR32X2TF \intadd_0/U2  ( .A(X_IN[7]), .B(DIVISION_HEAD[11]), .C(
        INTADD_0_N2), .CO(INTADD_0_N1), .S(\INTADD_0_SUM[6] ) );
  DFFRX2TF \rsht_bits_reg[3]  ( .D(N704), .CK(CLK), .RN(RST_N), .Q(
        \RSHT_BITS[3] ), .QN(N194) );
  DFFRX2TF \wtemp_reg[9]  ( .D(N673), .CK(CLK), .RN(RST_N), .Q(OPER_B[9]), 
        .QN(N193) );
  DFFRX2TF \wtemp_reg[12]  ( .D(N724), .CK(CLK), .RN(RST_N), .Q(OPER_B[12]), 
        .QN(N192) );
  DFFRX2TF \index_reg[3]  ( .D(N725), .CK(CLK), .RN(RST_N), .Q(N191), .QN(N124) );
  DFFRX2TF \wtemp_reg[11]  ( .D(N671), .CK(CLK), .RN(RST_N), .Q(OPER_B[11]), 
        .QN(N190) );
  DFFRX2TF \wtemp_reg[0]  ( .D(N682), .CK(CLK), .RN(RST_N), .Q(OPER_B[0]), 
        .QN(N189) );
  DFFRX2TF \wtemp_reg[3]  ( .D(N679), .CK(CLK), .RN(RST_N), .Q(OPER_B[3]), 
        .QN(N188) );
  DFFRX2TF \wtemp_reg[1]  ( .D(N681), .CK(CLK), .RN(RST_N), .Q(OPER_B[1]), 
        .QN(N187) );
  DFFRX2TF \index_reg[1]  ( .D(N699), .CK(CLK), .RN(RST_N), .Q(N186), .QN(N128) );
  DFFRX2TF \rsht_bits_reg[0]  ( .D(N703), .CK(CLK), .RN(RST_N), .Q(N185), .QN(
        N92) );
  DFFRX2TF \ytemp_reg[1]  ( .D(N693), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[1]), .QN(N184) );
  DFFRX2TF \ytemp_reg[0]  ( .D(N705), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[0]), .QN(N183) );
  DFFRX2TF sign_y_reg ( .D(N694), .CK(CLK), .RN(RST_N), .Q(SIGN_Y), .QN(N182)
         );
  DFFRX2TF \wtemp_reg[4]  ( .D(N678), .CK(CLK), .RN(RST_N), .Q(OPER_B[4]), 
        .QN(N181) );
  DFFSX2TF pre_work_reg ( .D(N695), .CK(CLK), .SN(RST_N), .Q(PRE_WORK), .QN(
        N180) );
  DFFRX2TF \xtemp_reg[12]  ( .D(N723), .CK(CLK), .RN(RST_N), .Q(XTEMP[12]), 
        .QN(N179) );
  DFFRX2TF \xtemp_reg[8]  ( .D(N711), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[12]), .QN(N178) );
  DFFRX2TF \ytemp_reg[6]  ( .D(N688), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[6]), .QN(N176) );
  DFFRX2TF \ytemp_reg[4]  ( .D(N690), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[4]), .QN(N175) );
  DFFRX2TF \ytemp_reg[10]  ( .D(N684), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[1]), .QN(N174) );
  DFFRX2TF \ytemp_reg[9]  ( .D(N685), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[0]), .QN(N173) );
  DFFRX2TF \ytemp_reg[7]  ( .D(N687), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[7]), .QN(N172) );
  DFFRX2TF \ytemp_reg[5]  ( .D(N689), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[5]), .QN(N171) );
  DFFRX2TF \ytemp_reg[3]  ( .D(N691), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[3]), .QN(N170) );
  DFFRX2TF \step_reg[0]  ( .D(N697), .CK(CLK), .RN(RST_N), .Q(N169), .QN(N122)
         );
  DFFRX2TF SEL_SRC_reg ( .D(N720), .CK(CLK), .RN(RST_N), .Q(POST_WORK), .QN(
        N168) );
  DFFRX2TF \ytemp_reg[11]  ( .D(N683), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[2]), .QN(N167) );
  DFFRX2TF \wtemp_reg[10]  ( .D(N672), .CK(CLK), .RN(RST_N), .Q(OPER_B[10]), 
        .QN(N166) );
  DFFRX2TF \wtemp_reg[8]  ( .D(N674), .CK(CLK), .RN(RST_N), .Q(OPER_B[8]), 
        .QN(N165) );
  DFFRX2TF \rsht_bits_reg[1]  ( .D(N702), .CK(CLK), .RN(RST_N), .Q(N164), .QN(
        N91) );
  DFFRX2TF \index_reg[0]  ( .D(N726), .CK(CLK), .RN(RST_N), .Q(N163), .QN(N129) );
  DFFRX2TF \wtemp_reg[2]  ( .D(N680), .CK(CLK), .RN(RST_N), .Q(OPER_B[2]), 
        .QN(N162) );
  DFFRX2TF \xtemp_reg[10]  ( .D(N709), .CK(CLK), .RN(RST_N), .Q(XTEMP[10]), 
        .QN(N161) );
  DFFRX2TF \xtemp_reg[6]  ( .D(N713), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[10]), .QN(N160) );
  DFFRX2TF \xtemp_reg[11]  ( .D(N708), .CK(CLK), .RN(RST_N), .Q(XTEMP[11]), 
        .QN(N159) );
  DFFRX2TF \xtemp_reg[5]  ( .D(N714), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[9]), .QN(N158) );
  DFFRX2TF \xtemp_reg[4]  ( .D(N715), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[8]), .QN(N157) );
  DFFRX2TF XOR_SRC_reg ( .D(N707), .CK(CLK), .RN(RST_N), .Q(N61), .QN(N73) );
  DFFRX2TF \xtemp_reg[0]  ( .D(N719), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[4]), .QN(N156) );
  DFFRX2TF \xtemp_reg[2]  ( .D(N717), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[6]), .QN(N155) );
  DFFRX2TF \xtemp_reg[7]  ( .D(N712), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[11]), .QN(N154) );
  DFFRX2TF \step_reg[3]  ( .D(N721), .CK(CLK), .RN(RST_N), .Q(STEP[3]), .QN(
        N153) );
  DFFRX2TF \step_reg[1]  ( .D(N700), .CK(CLK), .RN(RST_N), .Q(N152), .QN(N121)
         );
  DFFRX2TF \step_reg[2]  ( .D(N696), .CK(CLK), .RN(RST_N), .Q(STEP[2]), .QN(
        N151) );
  DFFRX2TF \ytemp_reg[2]  ( .D(N692), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[2]), .QN(N150) );
  DFFRX2TF \ytemp_reg[8]  ( .D(N686), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[8]), .QN(N149) );
  DFFRX2TF \rsht_bits_reg[2]  ( .D(N701), .CK(CLK), .RN(RST_N), .QN(N90) );
  DFFRX2TF SEL_Z_reg ( .D(N670), .CK(CLK), .RN(RST_N), .Q(N177), .QN(N123) );
  ADDHX1TF \add_x_132_1/U14  ( .A(OPER_B[0]), .B(OPER_A[0]), .CO(
        ADD_X_132_1_N13), .S(SUM_AB[0]) );
  CMPR32X2TF \add_x_132_1/U4  ( .A(OPER_A[10]), .B(OPER_B[10]), .C(
        ADD_X_132_1_N4), .CO(ADD_X_132_1_N3), .S(SUM_AB[10]) );
  CMPR32X2TF \add_x_132_1/U6  ( .A(OPER_A[8]), .B(OPER_B[8]), .C(
        ADD_X_132_1_N6), .CO(ADD_X_132_1_N5), .S(SUM_AB[8]) );
  CMPR32X2TF \add_x_132_1/U10  ( .A(OPER_A[4]), .B(OPER_B[4]), .C(
        ADD_X_132_1_N10), .CO(ADD_X_132_1_N9), .S(SUM_AB[4]) );
  CMPR32X2TF \add_x_132_1/U12  ( .A(OPER_A[2]), .B(OPER_B[2]), .C(
        ADD_X_132_1_N12), .CO(ADD_X_132_1_N11), .S(SUM_AB[2]) );
  CMPR32X2TF \add_x_132_1/U13  ( .A(OPER_A[1]), .B(OPER_B[1]), .C(
        ADD_X_132_1_N13), .CO(ADD_X_132_1_N12), .S(SUM_AB[1]) );
  CMPR32X2TF \add_x_132_1/U5  ( .A(OPER_A[9]), .B(OPER_B[9]), .C(
        ADD_X_132_1_N5), .CO(ADD_X_132_1_N4), .S(SUM_AB[9]) );
  CMPR32X2TF \add_x_132_1/U11  ( .A(OPER_A[3]), .B(OPER_B[3]), .C(
        ADD_X_132_1_N11), .CO(ADD_X_132_1_N10), .S(SUM_AB[3]) );
  CMPR32X2TF \add_x_132_1/U9  ( .A(OPER_A[5]), .B(OPER_B[5]), .C(
        ADD_X_132_1_N9), .CO(ADD_X_132_1_N8), .S(SUM_AB[5]) );
  CMPR32X2TF \add_x_132_1/U3  ( .A(OPER_A[11]), .B(OPER_B[11]), .C(
        ADD_X_132_1_N3), .CO(ADD_X_132_1_N2), .S(SUM_AB[11]) );
  DFFRX2TF sign_x_reg ( .D(N722), .CK(CLK), .RN(RST_N), .Q(N965), .QN(N74) );
  DFFRX1TF \ztemp_reg[0]  ( .D(N669), .CK(CLK), .RN(RST_N), .Q(ZTEMP[0]) );
  DFFRX1TF \wtemp_reg[6]  ( .D(N676), .CK(CLK), .RN(RST_N), .Q(OPER_B[6]) );
  DFFRX1TF \ztemp_reg[6]  ( .D(N663), .CK(CLK), .RN(RST_N), .Q(ZTEMP[6]) );
  DFFRX1TF \ztemp_reg[4]  ( .D(N665), .CK(CLK), .RN(RST_N), .Q(ZTEMP[4]) );
  DFFRX1TF \ztemp_reg[2]  ( .D(N667), .CK(CLK), .RN(RST_N), .Q(ZTEMP[2]) );
  DFFRX1TF \ztemp_reg[1]  ( .D(N668), .CK(CLK), .RN(RST_N), .Q(ZTEMP[1]) );
  DFFRX1TF \ztemp_reg[5]  ( .D(N664), .CK(CLK), .RN(RST_N), .Q(ZTEMP[5]) );
  DFFRX1TF \ztemp_reg[3]  ( .D(N666), .CK(CLK), .RN(RST_N), .Q(ZTEMP[3]) );
  DFFRX1TF \ztemp_reg[7]  ( .D(N662), .CK(CLK), .RN(RST_N), .Q(ZTEMP[7]) );
  DFFRX1TF \ztemp_reg[8]  ( .D(N661), .CK(CLK), .RN(RST_N), .Q(ZTEMP[8]) );
  DFFRX1TF \ztemp_reg[9]  ( .D(N660), .CK(CLK), .RN(RST_N), .Q(ZTEMP[9]) );
  DFFRX1TF \wtemp_reg[5]  ( .D(N677), .CK(CLK), .RN(RST_N), .Q(OPER_B[5]) );
  DFFRX1TF \wtemp_reg[7]  ( .D(N675), .CK(CLK), .RN(RST_N), .Q(OPER_B[7]) );
  DFFRX1TF \ztemp_reg[10]  ( .D(N659), .CK(CLK), .RN(RST_N), .Q(ZTEMP[10]) );
  DFFRX1TF \ztemp_reg[11]  ( .D(N658), .CK(CLK), .RN(RST_N), .Q(ZTEMP[11]) );
  DFFRX1TF \ztemp_reg[12]  ( .D(N657), .CK(CLK), .RN(RST_N), .Q(ZTEMP[12]) );
  DFFRX1TF \ytemp_reg[12]  ( .D(N706), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[3]), .QN(N649) );
  DFFRX2TF \xtemp_reg[1]  ( .D(N718), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[5]), .QN(N514) );
  DFFRX2TF \xtemp_reg[9]  ( .D(N710), .CK(CLK), .RN(RST_N), .Q(XTEMP[9]), .QN(
        N529) );
  DFFRX2TF \xtemp_reg[3]  ( .D(N716), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[7]), .QN(N423) );
  DFFRX2TF \index_reg[2]  ( .D(N698), .CK(CLK), .RN(RST_N), .Q(\INDEX[2] ) );
  NAND2X1TF U3 ( .A(N774), .B(N766), .Y(N394) );
  AOI222XLTF U4 ( .A0(DIVISION_HEAD[1]), .A1(DIVISION_HEAD[0]), .B0(
        DIVISION_HEAD[1]), .B1(N318), .C0(DIVISION_HEAD[0]), .C1(N317), .Y(
        N320) );
  NAND2X1TF U5 ( .A(ALU_START), .B(N263), .Y(N600) );
  OAI21X1TF U6 ( .A0(N893), .A1(N934), .B0(N932), .Y(N1) );
  AO21X1TF U7 ( .A0(N892), .A1(N937), .B0(N890), .Y(N2) );
  AOI22X1TF U8 ( .A0(OPER_A[7]), .A1(N1), .B0(OPER_B[7]), .B1(N2), .Y(N3) );
  OAI31X1TF U9 ( .A0(N892), .A1(N115), .A2(OPER_B[7]), .B0(N3), .Y(N4) );
  AOI211X1TF U10 ( .A0(C152_DATA4_7), .A1(N113), .B0(N211), .C0(N4), .Y(N5) );
  NAND3BX1TF U11 ( .AN(OPER_A[7]), .B(N893), .C(N931), .Y(N6) );
  OAI211X1TF U12 ( .A0(N894), .A1(N165), .B0(N5), .C0(N6), .Y(N675) );
  OAI211X1TF U13 ( .A0(N823), .A1(N376), .B0(N612), .C0(N640), .Y(N7) );
  AOI21XLTF U14 ( .A0(N377), .A1(N822), .B0(N7), .Y(N8) );
  NAND3X1TF U15 ( .A(N378), .B(N543), .C(N8), .Y(N9) );
  OAI22X1TF U16 ( .A0(N640), .A1(N764), .B0(N119), .B1(N379), .Y(N10) );
  OAI21X1TF U17 ( .A0(N10), .A1(N747), .B0(N9), .Y(N11) );
  OAI21X1TF U18 ( .A0(N168), .A1(N9), .B0(N11), .Y(N720) );
  AOI32X1TF U19 ( .A0(N116), .A1(N843), .A2(N935), .B0(N189), .B1(N843), .Y(
        N12) );
  AOI211X1TF U20 ( .A0(C152_DATA4_0), .A1(N114), .B0(N891), .C0(N12), .Y(N13)
         );
  OAI21X1TF U21 ( .A0(N854), .A1(N931), .B0(OPER_A[0]), .Y(N14) );
  OAI211X1TF U22 ( .A0(N187), .A1(N894), .B0(N13), .C0(N14), .Y(N682) );
  AOI22X1TF U23 ( .A0(N1011), .A1(ZTEMP[0]), .B0(N107), .B1(DIVISION_HEAD[0]), 
        .Y(N15) );
  AOI32XLTF U24 ( .A0(N1010), .A1(N15), .A2(N1019), .B0(N976), .B1(N15), .Y(
        N669) );
  OAI32X1TF U25 ( .A0(N190), .A1(N936), .A2(N116), .B0(N935), .B1(N190), .Y(
        N16) );
  CLKINVX1TF U26 ( .A(OPER_A[11]), .Y(N17) );
  OAI32X1TF U27 ( .A0(N17), .A1(N934), .A2(N933), .B0(N932), .B1(N17), .Y(N18)
         );
  AOI31X1TF U28 ( .A0(N933), .A1(N931), .A2(N17), .B0(N930), .Y(N19) );
  NOR2X1TF U29 ( .A(N115), .B(OPER_B[11]), .Y(N20) );
  AOI222XLTF U30 ( .A0(C152_DATA4_11), .A1(N113), .B0(N225), .B1(N964), .C0(
        N936), .C1(N20), .Y(N21) );
  OAI211X1TF U31 ( .A0(N192), .A1(N938), .B0(N19), .C0(N21), .Y(N22) );
  OR3X1TF U32 ( .A(N16), .B(N18), .C(N22), .Y(N671) );
  NOR2X1TF U33 ( .A(N933), .B(OPER_A[11]), .Y(N23) );
  XNOR2X1TF U34 ( .A(OPER_A[12]), .B(N23), .Y(N24) );
  AOI22X1TF U35 ( .A0(N24), .A1(N931), .B0(OPER_A[12]), .B1(N854), .Y(N25) );
  OAI21X1TF U36 ( .A0(N132), .A1(N549), .B0(N140), .Y(N26) );
  XNOR2X1TF U37 ( .A(N26), .B(N971), .Y(N27) );
  XNOR2X1TF U38 ( .A(DP_OP_333_124_4748_N1), .B(N27), .Y(N28) );
  NOR2X1TF U39 ( .A(OPER_B[11]), .B(N936), .Y(N29) );
  OAI31X1TF U40 ( .A0(N115), .A1(N29), .A2(OPER_B[12]), .B0(N825), .Y(N30) );
  AOI211X1TF U41 ( .A0(N114), .A1(N28), .B0(N930), .C0(N30), .Y(N31) );
  OAI31X1TF U42 ( .A0(OPER_B[11]), .A1(N936), .A2(N911), .B0(N874), .Y(N32) );
  AOI32X1TF U43 ( .A0(N130), .A1(OPER_B[12]), .A2(N32), .B0(N222), .B1(
        OPER_B[12]), .Y(N33) );
  NAND4BX1TF U44 ( .AN(N821), .B(N25), .C(N31), .D(N33), .Y(N724) );
  NOR3X1TF U45 ( .A(Y_IN[12]), .B(Y_IN[11]), .C(Y_IN[10]), .Y(N34) );
  NOR2X1TF U46 ( .A(N502), .B(N89), .Y(N35) );
  CLKINVX1TF U47 ( .A(Y_IN[6]), .Y(N36) );
  CLKINVX1TF U48 ( .A(N442), .Y(N37) );
  AOI22X1TF U49 ( .A0(N105), .A1(N738), .B0(N318), .B1(N37), .Y(N38) );
  OAI21X1TF U50 ( .A0(X_IN[4]), .A1(N317), .B0(N93), .Y(N39) );
  OAI22X1TF U51 ( .A0(N105), .A1(N738), .B0(X_IN[6]), .B1(N731), .Y(N40) );
  AOI31X1TF U52 ( .A0(N319), .A1(N38), .A2(N39), .B0(N40), .Y(N41) );
  AOI21X1TF U53 ( .A0(N731), .A1(X_IN[6]), .B0(N41), .Y(N42) );
  OA22X1TF U54 ( .A0(N43), .A1(N42), .B0(N488), .B1(N197), .Y(N44) );
  AO21X1TF U55 ( .A0(N468), .A1(N42), .B0(Y_IN[4]), .Y(N45) );
  AOI22X1TF U56 ( .A0(N488), .A1(N197), .B0(N44), .B1(N45), .Y(N46) );
  OA21XLTF U57 ( .A0(N36), .A1(N46), .B0(X_IN[9]), .Y(N47) );
  AOI211X1TF U58 ( .A0(N46), .A1(N36), .B0(N47), .C0(N35), .Y(N48) );
  AOI21X1TF U59 ( .A0(N502), .A1(Y_IN[7]), .B0(N48), .Y(N49) );
  AOI222XLTF U60 ( .A0(N762), .A1(N138), .B0(N762), .B1(N49), .C0(N138), .C1(
        N49), .Y(N50) );
  OAI21X1TF U61 ( .A0(Y_IN[9]), .A1(N305), .B0(N50), .Y(N51) );
  OAI211X1TF U62 ( .A0(X_IN[12]), .A1(N784), .B0(N34), .C0(N51), .Y(N770) );
  CLKINVX1TF U63 ( .A(X_IN[7]), .Y(N43) );
  NOR3X1TF U64 ( .A(N910), .B(N74), .C(N907), .Y(N52) );
  NOR2X1TF U65 ( .A(N166), .B(N938), .Y(N53) );
  AOI211X1TF U66 ( .A0(N113), .A1(C152_DATA4_9), .B0(N52), .C0(N53), .Y(N54)
         );
  NOR2X1TF U67 ( .A(N934), .B(OPER_A[9]), .Y(N55) );
  AOI22X1TF U68 ( .A0(SIGN_Y), .A1(N906), .B0(N909), .B1(N55), .Y(N56) );
  OAI21X1TF U69 ( .A0(N116), .A1(N908), .B0(N935), .Y(N57) );
  OAI21X1TF U70 ( .A0(N934), .A1(N909), .B0(N932), .Y(N58) );
  AOI22X1TF U71 ( .A0(OPER_B[9]), .A1(N57), .B0(OPER_A[9]), .B1(N58), .Y(N59)
         );
  NAND3X1TF U72 ( .A(N937), .B(N908), .C(N193), .Y(N60) );
  NAND4X1TF U73 ( .A(N54), .B(N56), .C(N59), .D(N60), .Y(N673) );
  INVX2TF U74 ( .A(N941), .Y(N118) );
  NOR3BX2TF U75 ( .AN(ALU_TYPE[2]), .B(ALU_TYPE[0]), .C(ALU_TYPE[1]), .Y(N263)
         );
  NOR3BXLTF U76 ( .AN(ALU_TYPE[0]), .B(ALU_TYPE[1]), .C(ALU_TYPE[2]), .Y(N262)
         );
  OAI32X4TF U77 ( .A0(N768), .A1(N767), .A2(X_IN[0]), .B0(N766), .B1(N768), 
        .Y(N771) );
  NOR2X4TF U78 ( .A(N385), .B(N769), .Y(N807) );
  OA21XLTF U79 ( .A0(SUM_AB[12]), .A1(N651), .B0(N119), .Y(N144) );
  NAND2X1TF U80 ( .A(N929), .B(N208), .Y(N221) );
  CLKINVX1TF U81 ( .A(SUM_AB[4]), .Y(N388) );
  AOI211X2TF U82 ( .A0(N571), .A1(N130), .B0(N595), .C0(N570), .Y(N597) );
  AO21X1TF U83 ( .A0(N777), .A1(N376), .B0(N823), .Y(N509) );
  CLKAND2X2TF U84 ( .A(N647), .B(N640), .Y(N546) );
  CLKINVX1TF U85 ( .A(N867), .Y(N865) );
  OR3X1TF U86 ( .A(PRE_WORK), .B(N606), .C(N600), .Y(N501) );
  AND2X2TF U87 ( .A(N117), .B(N195), .Y(N245) );
  CLKINVX1TF U88 ( .A(Y_IN[6]), .Y(N204) );
  AND2X2TF U89 ( .A(ZTEMP[0]), .B(N195), .Y(POUT[0]) );
  CLKINVX1TF U90 ( .A(N621), .Y(N623) );
  CLKINVX1TF U91 ( .A(N197), .Y(N205) );
  CLKINVX1TF U92 ( .A(N839), .Y(N834) );
  AOI211X1TF U93 ( .A0(N94), .A1(N747), .B0(N440), .C0(N439), .Y(N441) );
  AOI211X1TF U94 ( .A0(N106), .A1(N747), .B0(N458), .C0(N457), .Y(N459) );
  AOI211X1TF U95 ( .A0(N89), .A1(N747), .B0(N788), .C0(N787), .Y(N789) );
  OA21XLTF U96 ( .A0(SUM_AB[12]), .A1(N393), .B0(N119), .Y(N505) );
  AOI21X1TF U97 ( .A0(N767), .A1(N309), .B0(N385), .Y(N381) );
  CLKINVX2TF U98 ( .A(N871), .Y(N215) );
  INVX1TF U99 ( .A(N906), .Y(N889) );
  AND2X2TF U100 ( .A(N904), .B(N922), .Y(N937) );
  OAI21XLTF U101 ( .A0(N312), .A1(N629), .B0(N622), .Y(N313) );
  OR2X2TF U102 ( .A(N1011), .B(N133), .Y(N1012) );
  AOI22X1TF U103 ( .A0(Y_IN[9]), .A1(N802), .B0(X_IN[4]), .B1(N136), .Y(N803)
         );
  AOI21X1TF U104 ( .A0(N643), .A1(N130), .B0(N642), .Y(N646) );
  INVX1TF U105 ( .A(N403), .Y(N404) );
  OR2X2TF U106 ( .A(N385), .B(N764), .Y(N801) );
  OAI31XLTF U107 ( .A0(N119), .A1(N169), .A2(N632), .B0(N631), .Y(N637) );
  NAND3XLTF U108 ( .A(N130), .B(N824), .C(N823), .Y(N633) );
  AOI32XLTF U109 ( .A0(N822), .A1(N130), .A2(N823), .B0(N638), .B1(N130), .Y(
        N644) );
  OAI31X1TF U110 ( .A0(N565), .A1(N566), .A2(N564), .B0(N130), .Y(N582) );
  NAND4XLTF U111 ( .A(N612), .B(N611), .C(N610), .D(N609), .Y(N613) );
  OAI2BB2XLTF U112 ( .B0(N762), .B1(N804), .A0N(Y_IN[6]), .A1N(N802), .Y(N779)
         );
  INVX2TF U113 ( .A(N736), .Y(N99) );
  CLKINVX1TF U114 ( .A(OPER_A[1]), .Y(N832) );
  AOI22X1TF U115 ( .A0(DIVISION_HEAD[2]), .A1(N125), .B0(Y_IN[8]), .B1(N802), 
        .Y(N795) );
  INVX1TF U116 ( .A(OPER_A[0]), .Y(N831) );
  INVX1TF U117 ( .A(OPER_A[8]), .Y(N897) );
  INVX1TF U118 ( .A(OPER_A[6]), .Y(N881) );
  INVX1TF U119 ( .A(OPER_A[4]), .Y(N862) );
  AOI22X1TF U120 ( .A0(X_IN[2]), .A1(N802), .B0(N94), .B1(N444), .Y(N425) );
  INVX1TF U121 ( .A(OPER_A[10]), .Y(N915) );
  OAI211XLTF U122 ( .A0(N132), .A1(N368), .B0(N973), .C0(N601), .Y(N370) );
  AOI22X1TF U123 ( .A0(X_IN[2]), .A1(N444), .B0(X_IN[1]), .B1(N802), .Y(N417)
         );
  AOI22X1TF U124 ( .A0(Y_IN[1]), .A1(N802), .B0(DIVISION_REMA[4]), .B1(N125), 
        .Y(N732) );
  AOI22X1TF U125 ( .A0(N197), .A1(N802), .B0(N89), .B1(N791), .Y(N755) );
  NAND3BXLTF U126 ( .AN(N380), .B(N777), .C(N639), .Y(N369) );
  AOI22X1TF U127 ( .A0(XTEMP[10]), .A1(N95), .B0(X_IN[7]), .B1(N802), .Y(N480)
         );
  AOI22X1TF U128 ( .A0(Y_IN[3]), .A1(N802), .B0(DIVISION_REMA[6]), .B1(N125), 
        .Y(N742) );
  INVX2TF U129 ( .A(N132), .Y(N81) );
  AOI22X1TF U130 ( .A0(DIVISION_HEAD[2]), .A1(N110), .B0(ZTEMP[11]), .B1(N143), 
        .Y(N258) );
  AOI22X1TF U131 ( .A0(DIVISION_HEAD[3]), .A1(N110), .B0(ZTEMP[12]), .B1(N143), 
        .Y(N260) );
  AOI22X1TF U132 ( .A0(DIVISION_HEAD[1]), .A1(N110), .B0(ZTEMP[10]), .B1(N143), 
        .Y(N257) );
  INVX2TF U133 ( .A(N747), .Y(N97) );
  AOI22X1TF U134 ( .A0(DIVISION_REMA[0]), .A1(N109), .B0(ZTEMP[0]), .B1(N177), 
        .Y(N247) );
  AOI22X1TF U135 ( .A0(DIVISION_REMA[8]), .A1(N110), .B0(ZTEMP[8]), .B1(N177), 
        .Y(N255) );
  AOI22X1TF U136 ( .A0(DIVISION_REMA[7]), .A1(N110), .B0(ZTEMP[7]), .B1(N177), 
        .Y(N254) );
  AOI22X1TF U137 ( .A0(DIVISION_REMA[6]), .A1(N110), .B0(ZTEMP[6]), .B1(N177), 
        .Y(N253) );
  AOI22X1TF U138 ( .A0(DIVISION_REMA[5]), .A1(N110), .B0(ZTEMP[5]), .B1(N177), 
        .Y(N252) );
  AOI22X1TF U139 ( .A0(DIVISION_REMA[4]), .A1(N110), .B0(ZTEMP[4]), .B1(N177), 
        .Y(N251) );
  AND2X2TF U140 ( .A(N382), .B(N354), .Y(N736) );
  AOI22X1TF U141 ( .A0(DIVISION_REMA[3]), .A1(N110), .B0(ZTEMP[3]), .B1(N177), 
        .Y(N250) );
  AOI22X1TF U142 ( .A0(DIVISION_REMA[2]), .A1(N109), .B0(ZTEMP[2]), .B1(N177), 
        .Y(N249) );
  AOI22X1TF U143 ( .A0(DIVISION_HEAD[0]), .A1(N110), .B0(ZTEMP[9]), .B1(N143), 
        .Y(N256) );
  AOI22X1TF U144 ( .A0(DIVISION_REMA[1]), .A1(N109), .B0(ZTEMP[1]), .B1(N177), 
        .Y(N248) );
  OAI22X1TF U145 ( .A0(N133), .A1(N762), .B0(OFFSET[6]), .B1(N207), .Y(C2_Z_8)
         );
  INVX2TF U146 ( .A(N259), .Y(N109) );
  OAI22X1TF U147 ( .A0(N133), .A1(N805), .B0(OFFSET[9]), .B1(N140), .Y(C2_Z_11) );
  OAI22X1TF U148 ( .A0(N132), .A1(N548), .B0(OFFSET[8]), .B1(N140), .Y(C2_Z_10) );
  INVX2TF U149 ( .A(N813), .Y(N120) );
  OAI22X1TF U150 ( .A0(N133), .A1(N784), .B0(OFFSET[7]), .B1(N207), .Y(C2_Z_9)
         );
  OAI21XLTF U151 ( .A0(N132), .A1(N727), .B0(N207), .Y(C2_Z_0) );
  AND2X2TF U152 ( .A(N345), .B(N223), .Y(N941) );
  INVX1TF U153 ( .A(N345), .Y(N955) );
  AND2X2TF U154 ( .A(N354), .B(DP_OP_333_124_4748_N57), .Y(N747) );
  OR2X2TF U155 ( .A(N177), .B(N246), .Y(N259) );
  NAND2XLTF U156 ( .A(N223), .B(N946), .Y(N534) );
  AND2X2TF U157 ( .A(N123), .B(N246), .Y(N261) );
  OR2X2TF U158 ( .A(N351), .B(N600), .Y(N813) );
  CLKINVX2TF U159 ( .A(N500), .Y(N82) );
  AND2X2TF U160 ( .A(N224), .B(ALU_START), .Y(N971) );
  CLKAND2X2TF U161 ( .A(ZTEMP[11]), .B(N142), .Y(POUT[11]) );
  CLKAND2X2TF U162 ( .A(ZTEMP[7]), .B(N142), .Y(POUT[7]) );
  CLKAND2X2TF U163 ( .A(ZTEMP[6]), .B(N142), .Y(POUT[6]) );
  CLKAND2X2TF U164 ( .A(ZTEMP[10]), .B(N142), .Y(POUT[10]) );
  CLKAND2X2TF U165 ( .A(ZTEMP[9]), .B(N142), .Y(POUT[9]) );
  CLKAND2X2TF U166 ( .A(ZTEMP[8]), .B(N142), .Y(POUT[8]) );
  AOI22X1TF U167 ( .A0(N73), .A1(DIVISION_HEAD[3]), .B0(XTEMP[12]), .B1(N61), 
        .Y(N349) );
  INVX2TF U168 ( .A(N73), .Y(N117) );
  CLKAND2X2TF U169 ( .A(ZTEMP[12]), .B(N195), .Y(POUT[12]) );
  CLKAND2X2TF U170 ( .A(ZTEMP[2]), .B(N195), .Y(POUT[2]) );
  CLKAND2X2TF U171 ( .A(ZTEMP[4]), .B(N195), .Y(POUT[4]) );
  CLKAND2X2TF U172 ( .A(ZTEMP[1]), .B(N195), .Y(POUT[1]) );
  INVX2TF U173 ( .A(N198), .Y(N89) );
  CLKAND2X2TF U174 ( .A(ZTEMP[3]), .B(N195), .Y(POUT[3]) );
  AND2X2TF U175 ( .A(N195), .B(N73), .Y(N244) );
  INVX2TF U176 ( .A(N200), .Y(N105) );
  AND2X1TF U177 ( .A(\INDEX[2] ), .B(N625), .Y(N314) );
  CLKAND2X2TF U178 ( .A(ZTEMP[5]), .B(N195), .Y(POUT[5]) );
  NAND2XLTF U179 ( .A(DIVISION_HEAD[4]), .B(N263), .Y(N226) );
  INVX2TF U180 ( .A(X_IN[3]), .Y(N199) );
  INVX2TF U181 ( .A(X_IN[5]), .Y(N200) );
  INVX2TF U182 ( .A(ALU_TYPE[1]), .Y(N202) );
  INVX2TF U183 ( .A(X_IN[11]), .Y(N201) );
  INVX2TF U184 ( .A(Y_IN[7]), .Y(N198) );
  INVX2TF U185 ( .A(N244), .Y(N83) );
  INVX2TF U186 ( .A(N244), .Y(N84) );
  INVX2TF U187 ( .A(N245), .Y(N85) );
  INVX2TF U188 ( .A(N245), .Y(N86) );
  INVX2TF U189 ( .A(N1019), .Y(N87) );
  INVX2TF U190 ( .A(N1019), .Y(N88) );
  INVX2TF U191 ( .A(N199), .Y(N93) );
  INVX2TF U192 ( .A(N199), .Y(N94) );
  INVX2TF U193 ( .A(N501), .Y(N95) );
  INVX2TF U194 ( .A(N501), .Y(N96) );
  INVX2TF U195 ( .A(N747), .Y(N98) );
  INVX2TF U196 ( .A(N736), .Y(N100) );
  INVX2TF U197 ( .A(N394), .Y(N101) );
  INVX2TF U198 ( .A(N394), .Y(N102) );
  INVX2TF U199 ( .A(N263), .Y(N103) );
  INVX2TF U200 ( .A(N263), .Y(N104) );
  INVX2TF U201 ( .A(N200), .Y(N106) );
  INVX2TF U202 ( .A(N1012), .Y(N107) );
  INVX2TF U203 ( .A(N1012), .Y(N108) );
  INVX2TF U204 ( .A(N259), .Y(N110) );
  INVX2TF U205 ( .A(N261), .Y(N111) );
  INVX2TF U206 ( .A(N261), .Y(N112) );
  INVX2TF U207 ( .A(N221), .Y(N113) );
  INVX2TF U208 ( .A(N221), .Y(N114) );
  INVX2TF U209 ( .A(N937), .Y(N115) );
  INVX2TF U210 ( .A(N937), .Y(N116) );
  INVX2TF U211 ( .A(N941), .Y(N119) );
  INVX2TF U212 ( .A(N813), .Y(N125) );
  INVX2TF U213 ( .A(N509), .Y(N126) );
  INVX2TF U214 ( .A(N509), .Y(N127) );
  INVX2TF U215 ( .A(N118), .Y(N130) );
  INVX2TF U216 ( .A(N99), .Y(N131) );
  INVX2TF U217 ( .A(N971), .Y(N132) );
  INVX2TF U218 ( .A(N971), .Y(N133) );
  AOI222X4TF U219 ( .A0(N487), .A1(N161), .B0(N487), .B1(N502), .C0(N161), 
        .C1(N502), .Y(N497) );
  NOR2X2TF U220 ( .A(N342), .B(N956), .Y(N354) );
  NOR3X2TF U221 ( .A(N118), .B(N605), .C(N632), .Y(N618) );
  INVX2TF U222 ( .A(N505), .Y(N134) );
  INVX2TF U223 ( .A(N505), .Y(N135) );
  INVX2TF U224 ( .A(N801), .Y(N136) );
  INVX2TF U225 ( .A(N801), .Y(N137) );
  NAND2X2TF U226 ( .A(N123), .B(N763), .Y(N454) );
  AOI21X2TF U227 ( .A0(N941), .A1(N921), .B0(N222), .Y(N935) );
  INVX2TF U228 ( .A(N201), .Y(N138) );
  INVX2TF U229 ( .A(N201), .Y(N139) );
  AOI211XLTF U230 ( .A0(N832), .A1(N831), .B0(OPER_A[2]), .C0(N916), .Y(N833)
         );
  OAI32XLTF U231 ( .A0(OPER_A[8]), .A1(N898), .A2(N916), .B0(N897), .B1(N896), 
        .Y(N899) );
  OAI32XLTF U232 ( .A0(OPER_A[10]), .A1(N917), .A2(N916), .B0(N915), .B1(N914), 
        .Y(N918) );
  OAI32XLTF U233 ( .A0(OPER_A[6]), .A1(N882), .A2(N916), .B0(N881), .B1(N880), 
        .Y(N883) );
  INVXLTF U234 ( .A(N916), .Y(N913) );
  INVXLTF U235 ( .A(X_IN[2]), .Y(N772) );
  INVX2TF U236 ( .A(DP_OP_333_124_4748_N57), .Y(N140) );
  INVX2TF U237 ( .A(N969), .Y(N141) );
  AOI2BB1X2TF U238 ( .A0N(N963), .A1N(N962), .B0(N961), .Y(N1011) );
  CLKBUFX2TF U239 ( .A(N195), .Y(N142) );
  CLKBUFX2TF U240 ( .A(N262), .Y(N195) );
  NOR3XLTF U241 ( .A(N73), .B(N910), .C(N972), .Y(N821) );
  NAND2X2TF U242 ( .A(N970), .B(N929), .Y(N910) );
  AOI21XLTF U243 ( .A0(N824), .A1(N823), .B0(N822), .Y(N835) );
  INVXLTF U244 ( .A(N822), .Y(N379) );
  NOR3BX4TF U245 ( .AN(N384), .B(N381), .C(N131), .Y(N513) );
  AOI222X4TF U246 ( .A0(XTEMP[9]), .A1(X_IN[9]), .B0(XTEMP[9]), .B1(N478), 
        .C0(X_IN[9]), .C1(N478), .Y(N487) );
  AOI222X4TF U247 ( .A0(N178), .A1(N488), .B0(N178), .B1(N464), .C0(N488), 
        .C1(N464), .Y(N478) );
  OAI31XLTF U248 ( .A0(OPER_A[1]), .A1(N916), .A2(OPER_A[0]), .B0(N837), .Y(
        N838) );
  OAI21X2TF U249 ( .A0(N514), .A1(N111), .B0(N248), .Y(OPER_A[1]) );
  INVX2TF U250 ( .A(N123), .Y(N143) );
  NAND2X2TF U251 ( .A(N763), .B(N143), .Y(N559) );
  AOI22XLTF U252 ( .A0(X_IN[1]), .A1(N807), .B0(X_IN[0]), .B1(N136), .Y(N754)
         );
  AOI22XLTF U253 ( .A0(X_IN[4]), .A1(N101), .B0(X_IN[6]), .B1(N807), .Y(N552)
         );
  AOI22XLTF U254 ( .A0(X_IN[12]), .A1(N807), .B0(N139), .B1(N136), .Y(N436) );
  AOI22XLTF U255 ( .A0(X_IN[2]), .A1(N101), .B0(X_IN[4]), .B1(N807), .Y(N792)
         );
  AOI22XLTF U256 ( .A0(DIVISION_HEAD[5]), .A1(N95), .B0(X_IN[7]), .B1(N807), 
        .Y(N387) );
  AOI22XLTF U257 ( .A0(X_IN[10]), .A1(N136), .B0(N139), .B1(N807), .Y(N427) );
  AOI22XLTF U258 ( .A0(X_IN[2]), .A1(N136), .B0(N94), .B1(N807), .Y(N786) );
  AOI22XLTF U259 ( .A0(N94), .A1(N101), .B0(N106), .B1(N807), .Y(N808) );
  NAND2X2TF U260 ( .A(PRE_WORK), .B(N971), .Y(N385) );
  NOR4X2TF U261 ( .A(N648), .B(N943), .C(N370), .D(N369), .Y(N642) );
  NOR2X2TF U262 ( .A(N342), .B(N604), .Y(N566) );
  NOR2BX2TF U263 ( .AN(N544), .B(N382), .Y(N629) );
  NOR2X2TF U264 ( .A(N351), .B(N132), .Y(N382) );
  INVX2TF U265 ( .A(N144), .Y(N145) );
  INVX2TF U266 ( .A(N144), .Y(N146) );
  AOI22X2TF U267 ( .A0(N349), .A1(N347), .B0(N940), .B1(N350), .Y(N922) );
  NOR3X4TF U268 ( .A(N202), .B(ALU_TYPE[0]), .C(ALU_TYPE[2]), .Y(N224) );
  XNOR2X1TF U269 ( .A(OPER_A[12]), .B(ADD_X_132_1_N2), .Y(N147) );
  CMPR32X2TF U270 ( .A(OPER_A[7]), .B(OPER_B[7]), .C(ADD_X_132_1_N7), .CO(
        ADD_X_132_1_N6), .S(SUM_AB[7]) );
  CMPR32X2TF U271 ( .A(OPER_A[6]), .B(OPER_B[6]), .C(ADD_X_132_1_N8), .CO(
        ADD_X_132_1_N7), .S(SUM_AB[6]) );
  XNOR2X2TF U272 ( .A(N147), .B(OPER_B[12]), .Y(SUM_AB[12]) );
  AOI32X1TF U273 ( .A0(N941), .A1(N61), .A2(N564), .B0(N618), .B1(N73), .Y(
        N545) );
  AOI22X1TF U274 ( .A0(N73), .A1(N168), .B0(POST_WORK), .B1(N117), .Y(N246) );
  OAI31X1TF U275 ( .A0(N133), .A1(N949), .A2(N948), .B0(N947), .Y(N950) );
  NAND2X1TF U276 ( .A(N317), .B(N727), .Y(N319) );
  NAND2X1TF U277 ( .A(N477), .B(N476), .Y(N486) );
  NOR2X1TF U278 ( .A(SUM_AB[8]), .B(N462), .Y(N477) );
  OA22X1TF U279 ( .A0(N769), .A1(N558), .B0(N764), .B1(N765), .Y(N309) );
  INVX2TF U280 ( .A(N929), .Y(N222) );
  OAI21X1TF U281 ( .A0(N948), .A1(N610), .B0(N647), .Y(N961) );
  NAND2X1TF U282 ( .A(Y_IN[1]), .B(Y_IN[0]), .Y(N318) );
  NOR2X1TF U283 ( .A(SUM_AB[10]), .B(N486), .Y(N499) );
  NOR2X2TF U284 ( .A(N222), .B(N118), .Y(N904) );
  OR2X2TF U285 ( .A(N961), .B(N203), .Y(N929) );
  NOR2X1TF U286 ( .A(\INDEX[2] ), .B(N621), .Y(N312) );
  NAND2X1TF U287 ( .A(N129), .B(N128), .Y(N621) );
  OAI21X1TF U288 ( .A0(DIVISION_HEAD[12]), .A1(N549), .B0(N341), .Y(N948) );
  AOI2BB1X1TF U289 ( .A0N(DIVISION_HEAD[6]), .A1N(N330), .B0(Y_IN[6]), .Y(N328) );
  AOI21X1TF U290 ( .A0(N197), .A1(N514), .B0(N327), .Y(N330) );
  AOI2BB1X1TF U291 ( .A0N(DIVISION_HEAD[4]), .A1N(N326), .B0(Y_IN[4]), .Y(N324) );
  NOR2X1TF U292 ( .A(Y_IN[3]), .B(N649), .Y(N322) );
  AOI211X1TF U293 ( .A0(Y_IN[11]), .A1(N305), .B0(Y_IN[12]), .C0(N287), .Y(
        N767) );
  NAND2X1TF U294 ( .A(N912), .B(N904), .Y(N932) );
  NAND2X1TF U295 ( .A(N565), .B(N350), .Y(N916) );
  AOI2BB1X1TF U296 ( .A0N(N608), .A1N(N346), .B0(N962), .Y(N203) );
  NOR2X1TF U297 ( .A(PRE_WORK), .B(N343), .Y(N345) );
  NAND2X1TF U298 ( .A(N122), .B(N152), .Y(N605) );
  NOR2X1TF U299 ( .A(N124), .B(N628), .Y(N343) );
  NAND2X1TF U300 ( .A(N566), .B(N382), .Y(N610) );
  NAND2X1TF U301 ( .A(N180), .B(N368), .Y(N351) );
  NAND2X1TF U302 ( .A(N151), .B(N153), .Y(N342) );
  NAND2X1TF U303 ( .A(N454), .B(N460), .Y(N471) );
  NAND2X2TF U304 ( .A(N547), .B(N384), .Y(N460) );
  CLKBUFX2TF U305 ( .A(N782), .Y(N196) );
  NAND2X1TF U306 ( .A(N121), .B(N122), .Y(N956) );
  NAND3X1TF U307 ( .A(N962), .B(N132), .C(N600), .Y(N647) );
  AND2X2TF U308 ( .A(ALU_START), .B(N142), .Y(N223) );
  NAND2X1TF U309 ( .A(N124), .B(N312), .Y(N368) );
  NAND2X1TF U310 ( .A(N121), .B(N169), .Y(N604) );
  CLKBUFX2TF U311 ( .A(Y_IN[5]), .Y(N197) );
  NOR3X1TF U312 ( .A(N606), .B(N605), .C(N777), .Y(N607) );
  OR3X1TF U313 ( .A(N888), .B(N887), .C(N217), .Y(N676) );
  OAI2BB2XLTF U314 ( .B0(N889), .B1(N972), .A0N(C152_DATA4_6), .A1N(N113), .Y(
        N217) );
  OAI2BB2XLTF U315 ( .B0(N886), .B1(N924), .A0N(N222), .A1N(OPER_B[6]), .Y(
        N887) );
  INVX2TF U316 ( .A(N460), .Y(N475) );
  AOI32X1TF U317 ( .A0(N970), .A1(N969), .A2(N968), .B0(N130), .B1(N969), .Y(
        N1019) );
  NAND2X1TF U318 ( .A(N647), .B(N97), .Y(N944) );
  NAND2X1TF U319 ( .A(N566), .B(DP_OP_333_124_4748_N57), .Y(N393) );
  NAND2X1TF U320 ( .A(N960), .B(DP_OP_333_124_4748_N57), .Y(N651) );
  INVX2TF U321 ( .A(N367), .Y(N763) );
  NAND2X1TF U322 ( .A(N382), .B(N960), .Y(N367) );
  NOR2BX2TF U323 ( .AN(N547), .B(N557), .Y(N814) );
  NOR2X1TF U324 ( .A(N180), .B(N600), .Y(N356) );
  NAND2X1TF U325 ( .A(SIGN_Y), .B(N965), .Y(N972) );
  NAND2X1TF U326 ( .A(N904), .B(N877), .Y(N894) );
  INVX2TF U327 ( .A(DP_OP_333_124_4748_N57), .Y(N207) );
  AND2X2TF U328 ( .A(N223), .B(PRE_WORK), .Y(DP_OP_333_124_4748_N57) );
  AOI21X1TF U329 ( .A0(N949), .A1(N967), .B0(N366), .Y(N970) );
  NAND2X1TF U330 ( .A(N151), .B(STEP[3]), .Y(N632) );
  NOR2X2TF U331 ( .A(N342), .B(N605), .Y(N960) );
  INVX2TF U332 ( .A(N223), .Y(N962) );
  AO22X1TF U333 ( .A0(N375), .A1(XTEMP[12]), .B0(N363), .B1(N965), .Y(N722) );
  AOI211X1TF U334 ( .A0(N223), .A1(N608), .B0(N945), .C0(N607), .Y(N611) );
  AOI32X1TF U335 ( .A0(N967), .A1(N364), .A2(N958), .B0(N973), .B1(N364), .Y(
        N365) );
  NAND2X1TF U336 ( .A(N643), .B(N125), .Y(N615) );
  NAND2X1TF U337 ( .A(N946), .B(DP_OP_333_124_4748_N57), .Y(N635) );
  NAND2X1TF U338 ( .A(N114), .B(C152_DATA4_8), .Y(N218) );
  OAI22X1TF U339 ( .A0(N514), .A1(N99), .B0(N155), .B1(N454), .Y(N405) );
  AOI32X1TF U340 ( .A0(N126), .A1(DIVISION_HEAD[4]), .A2(N750), .B0(N471), 
        .B1(DIVISION_HEAD[4]), .Y(N391) );
  OAI22X1TF U341 ( .A0(N529), .A1(N100), .B0(N488), .B1(N98), .Y(N489) );
  INVX2TF U342 ( .A(N1015), .Y(N1010) );
  OAI2BB2XLTF U343 ( .B0(N61), .B1(N972), .A0N(N972), .A1N(N61), .Y(N974) );
  OAI22X1TF U344 ( .A0(N161), .A1(N99), .B0(N500), .B1(N97), .Y(N504) );
  INVX2TF U345 ( .A(N120), .Y(N777) );
  NOR2X2TF U346 ( .A(N763), .B(N196), .Y(N761) );
  NAND2X1TF U347 ( .A(N354), .B(N120), .Y(N544) );
  NAND2X1TF U348 ( .A(N132), .B(N140), .Y(N208) );
  NOR2X1TF U349 ( .A(N956), .B(N632), .Y(N564) );
  OAI21X2TF U350 ( .A0(N156), .A1(N111), .B0(N247), .Y(OPER_A[0]) );
  NOR2X1TF U351 ( .A(N605), .B(N954), .Y(N565) );
  NAND2X1TF U352 ( .A(STEP[2]), .B(N153), .Y(N954) );
  OAI32X1TF U353 ( .A0(N650), .A1(N182), .A2(N944), .B0(N649), .B1(N651), .Y(
        N694) );
  OAI21X1TF U354 ( .A0(N180), .A1(N648), .B0(N647), .Y(N695) );
  AOI22X1TF U355 ( .A0(N543), .A1(N73), .B0(N542), .B1(N541), .Y(N707) );
  INVX2TF U356 ( .A(N543), .Y(N541) );
  OAI31X1TF U357 ( .A0(N540), .A1(N539), .A2(N538), .B0(N537), .Y(N542) );
  AOI211X1TF U358 ( .A0(N536), .A1(XTEMP[12]), .B0(N535), .C0(N534), .Y(N537)
         );
  OAI31X1TF U359 ( .A0(DIVISION_HEAD[1]), .A1(N533), .A2(N161), .B0(N532), .Y(
        N536) );
  AOI22X1TF U360 ( .A0(N531), .A1(N530), .B0(XTEMP[11]), .B1(N167), .Y(N532)
         );
  OAI22X1TF U361 ( .A0(DIVISION_HEAD[0]), .A1(N529), .B0(DIVISION_REMA[8]), 
        .B1(N178), .Y(N530) );
  INVX2TF U362 ( .A(N539), .Y(N531) );
  NOR2X1TF U363 ( .A(XTEMP[11]), .B(N167), .Y(N533) );
  OAI22X1TF U364 ( .A0(DIVISION_HEAD[12]), .A1(N149), .B0(XTEMP[12]), .B1(N649), .Y(N538) );
  OAI21X1TF U365 ( .A0(XTEMP[11]), .A1(N167), .B0(N528), .Y(N539) );
  AOI22X1TF U366 ( .A0(DIVISION_HEAD[0]), .A1(N529), .B0(DIVISION_HEAD[1]), 
        .B1(N161), .Y(N528) );
  AOI21X1TF U367 ( .A0(DIVISION_HEAD[11]), .A1(N172), .B0(N527), .Y(N540) );
  AOI211X1TF U368 ( .A0(DIVISION_REMA[6]), .A1(N160), .B0(N526), .C0(N525), 
        .Y(N527) );
  NOR2X1TF U369 ( .A(DIVISION_HEAD[11]), .B(N172), .Y(N525) );
  AOI21X1TF U370 ( .A0(DIVISION_HEAD[9]), .A1(N171), .B0(N523), .Y(N524) );
  AOI211X1TF U371 ( .A0(DIVISION_REMA[4]), .A1(N157), .B0(N522), .C0(N521), 
        .Y(N523) );
  NOR2X1TF U372 ( .A(DIVISION_HEAD[9]), .B(N171), .Y(N521) );
  AOI21X1TF U373 ( .A0(DIVISION_HEAD[7]), .A1(N170), .B0(N519), .Y(N520) );
  AOI211X1TF U374 ( .A0(N518), .A1(DIVISION_REMA[2]), .B0(N517), .C0(N516), 
        .Y(N519) );
  NOR2X1TF U375 ( .A(DIVISION_HEAD[7]), .B(N170), .Y(N517) );
  OAI21X1TF U376 ( .A0(DIVISION_HEAD[5]), .A1(N184), .B0(N515), .Y(N518) );
  OAI211X1TF U377 ( .A0(DIVISION_REMA[1]), .A1(N514), .B0(DIVISION_REMA[0]), 
        .C0(N156), .Y(N515) );
  OAI21X1TF U378 ( .A0(N123), .A1(N952), .B0(N951), .Y(N670) );
  OAI21X1TF U379 ( .A0(N950), .A1(N970), .B0(N952), .Y(N951) );
  OR4X2TF U380 ( .A(N945), .B(N944), .C(N943), .D(N942), .Y(N952) );
  OAI22X1TF U381 ( .A0(N119), .A1(N940), .B0(N939), .B1(N973), .Y(N942) );
  OAI21X1TF U382 ( .A0(N597), .A1(N586), .B0(N585), .Y(N702) );
  AOI31X1TF U383 ( .A0(N584), .A1(N589), .A2(N591), .B0(N583), .Y(N586) );
  OAI22X1TF U384 ( .A0(N128), .A1(N582), .B0(N593), .B1(N589), .Y(N583) );
  OAI21X1TF U385 ( .A0(N128), .A1(N620), .B0(N619), .Y(N699) );
  AOI31X1TF U386 ( .A0(N618), .A1(N621), .A2(N617), .B0(N616), .Y(N619) );
  OAI32X1TF U387 ( .A0(N629), .A1(N630), .A2(N621), .B0(N617), .B1(N629), .Y(
        N616) );
  AOI22X1TF U388 ( .A0(N597), .A1(N92), .B0(N581), .B1(N580), .Y(N703) );
  AOI211X1TF U389 ( .A0(N595), .A1(N163), .B0(N579), .C0(N791), .Y(N581) );
  AOI21X1TF U390 ( .A0(N578), .A1(N777), .B0(N185), .Y(N579) );
  OAI31X1TF U391 ( .A0(N630), .A1(N629), .A2(N628), .B0(N627), .Y(N698) );
  AOI22X1TF U392 ( .A0(\INDEX[2] ), .A1(N626), .B0(N625), .B1(N624), .Y(N627)
         );
  OAI21X1TF U393 ( .A0(N623), .A1(N629), .B0(N622), .Y(N626) );
  OAI211X1TF U394 ( .A0(N119), .A1(N372), .B0(N645), .C0(N371), .Y(N721) );
  AOI22X1TF U395 ( .A0(STEP[3]), .A1(N642), .B0(N377), .B1(N574), .Y(N371) );
  OAI211X1TF U396 ( .A0(N183), .A1(N615), .B0(N631), .C0(N614), .Y(N700) );
  AOI21X1TF U397 ( .A0(N642), .A1(N152), .B0(N613), .Y(N614) );
  NOR3X1TF U398 ( .A(STEP[3]), .B(N119), .C(N604), .Y(N945) );
  AOI211X1TF U399 ( .A0(N824), .A1(N377), .B0(N375), .C0(N374), .Y(N612) );
  AOI21X1TF U400 ( .A0(N383), .A1(N373), .B0(N777), .Y(N374) );
  NOR2X1TF U401 ( .A(N118), .B(N823), .Y(N377) );
  OAI22X1TF U402 ( .A0(N90), .A1(N598), .B0(N597), .B1(N596), .Y(N701) );
  AOI21X1TF U403 ( .A0(\INDEX[2] ), .A1(N595), .B0(N594), .Y(N596) );
  OAI22X1TF U404 ( .A0(N593), .A1(N592), .B0(N591), .B1(N590), .Y(N594) );
  INVX2TF U405 ( .A(N588), .Y(N593) );
  AOI21X1TF U406 ( .A0(N589), .A1(N588), .B0(N587), .Y(N598) );
  OAI211X1TF U407 ( .A0(N646), .A1(N151), .B0(N645), .C0(N644), .Y(N696) );
  NOR2X1TF U408 ( .A(N650), .B(N365), .Y(N645) );
  INVX2TF U409 ( .A(N651), .Y(N650) );
  OAI22X1TF U410 ( .A0(N169), .A1(N954), .B0(N823), .B1(N967), .Y(N638) );
  AOI211X1TF U411 ( .A0(N642), .A1(N169), .B0(N637), .C0(N636), .Y(N641) );
  AOI21X1TF U412 ( .A0(N81), .A1(N603), .B0(N602), .Y(N631) );
  OAI21X1TF U413 ( .A0(N601), .A1(N600), .B0(N599), .Y(N602) );
  OAI22X1TF U414 ( .A0(N597), .A1(N577), .B0(N576), .B1(N194), .Y(N704) );
  AOI21X1TF U415 ( .A0(N592), .A1(N588), .B0(N587), .Y(N576) );
  OAI21X1TF U416 ( .A0(N90), .A1(N591), .B0(N584), .Y(N590) );
  INVX2TF U417 ( .A(N615), .Y(N584) );
  INVX2TF U418 ( .A(N597), .Y(N580) );
  OAI31X1TF U419 ( .A0(N606), .A1(N605), .A2(N777), .B0(N578), .Y(N588) );
  OAI32X1TF U420 ( .A0(N575), .A1(N824), .A2(N574), .B0(N130), .B1(N575), .Y(
        N578) );
  INVX2TF U421 ( .A(N573), .Y(N575) );
  AOI21X1TF U422 ( .A0(N595), .A1(N191), .B0(N572), .Y(N577) );
  AOI32X1TF U423 ( .A0(N566), .A1(N125), .A2(N183), .B0(N960), .B1(N120), .Y(
        N568) );
  AOI31X1TF U424 ( .A0(N130), .A1(N824), .A2(N823), .B0(N944), .Y(N569) );
  INVX2TF U425 ( .A(N582), .Y(N595) );
  AOI32X1TF U426 ( .A0(N314), .A1(N124), .A2(N618), .B0(N191), .B1(N313), .Y(
        N316) );
  NOR2X1TF U427 ( .A(N630), .B(N624), .Y(N622) );
  AOI21X1TF U428 ( .A0(\INDEX[2] ), .A1(N625), .B0(N378), .Y(N624) );
  INVX2TF U429 ( .A(N620), .Y(N630) );
  INVX2TF U430 ( .A(N617), .Y(N625) );
  OAI21X1TF U431 ( .A0(N129), .A1(N620), .B0(N311), .Y(N726) );
  OAI21X1TF U432 ( .A0(N310), .A1(N381), .B0(N620), .Y(N311) );
  AOI32X1TF U433 ( .A0(N629), .A1(N635), .A2(N378), .B0(N163), .B1(N635), .Y(
        N310) );
  INVX2TF U434 ( .A(N265), .Y(N634) );
  AOI31X1TF U435 ( .A0(N956), .A1(N373), .A2(N383), .B0(N777), .Y(N265) );
  OAI21X1TF U436 ( .A0(N354), .A1(N264), .B0(N941), .Y(N364) );
  AOI22X1TF U437 ( .A0(N903), .A1(N904), .B0(N222), .B1(OPER_B[8]), .Y(N219)
         );
  OAI21X1TF U438 ( .A0(N902), .A1(N165), .B0(N901), .Y(N903) );
  AOI211X1TF U439 ( .A0(N920), .A1(OPER_B[9]), .B0(N900), .C0(N899), .Y(N901)
         );
  AOI21X1TF U440 ( .A0(N913), .A1(N898), .B0(N912), .Y(N896) );
  NOR3X1TF U441 ( .A(N911), .B(OPER_B[8]), .C(N895), .Y(N900) );
  AOI21X1TF U442 ( .A0(N895), .A1(N922), .B0(N921), .Y(N902) );
  OAI21X1TF U443 ( .A0(N450), .A1(N449), .B0(N460), .Y(N451) );
  AOI22X1TF U444 ( .A0(DIVISION_HEAD[11]), .A1(N96), .B0(X_IN[12]), .B1(N137), 
        .Y(N445) );
  AOI22X1TF U445 ( .A0(N106), .A1(N444), .B0(N139), .B1(N102), .Y(N446) );
  AOI22X1TF U446 ( .A0(SUM_AB[6]), .A1(N134), .B0(N493), .B1(N992), .Y(N447)
         );
  OAI22X1TF U447 ( .A0(N158), .A1(N100), .B0(N442), .B1(N98), .Y(N450) );
  INVX2TF U448 ( .A(N888), .Y(N214) );
  AOI31X1TF U449 ( .A0(N842), .A1(N841), .A2(N840), .B0(N924), .Y(N844) );
  AOI32X1TF U450 ( .A0(N839), .A1(OPER_B[2]), .A2(N922), .B0(N921), .B1(
        OPER_B[2]), .Y(N840) );
  AOI22X1TF U451 ( .A0(N920), .A1(OPER_B[3]), .B0(OPER_A[2]), .B1(N838), .Y(
        N841) );
  AOI31X1TF U452 ( .A0(N922), .A1(N162), .A2(N834), .B0(N833), .Y(N842) );
  OAI211X1TF U453 ( .A0(N1010), .A1(N985), .B0(N984), .C0(N983), .Y(N666) );
  AOI22X1TF U454 ( .A0(DIVISION_HEAD[3]), .A1(N107), .B0(ZTEMP[3]), .B1(N1011), 
        .Y(N984) );
  OAI211X1TF U455 ( .A0(N1010), .A1(N991), .B0(N990), .C0(N989), .Y(N664) );
  AOI22X1TF U456 ( .A0(DIVISION_HEAD[5]), .A1(N107), .B0(ZTEMP[5]), .B1(N141), 
        .Y(N990) );
  OAI211X1TF U457 ( .A0(N1010), .A1(N1003), .B0(N1002), .C0(N1001), .Y(N660)
         );
  AOI22X1TF U458 ( .A0(DIVISION_HEAD[9]), .A1(N107), .B0(ZTEMP[9]), .B1(N1011), 
        .Y(N1002) );
  OAI211X1TF U459 ( .A0(N1010), .A1(N997), .B0(N996), .C0(N995), .Y(N662) );
  AOI22X1TF U460 ( .A0(DIVISION_HEAD[7]), .A1(N107), .B0(ZTEMP[7]), .B1(N141), 
        .Y(N996) );
  AOI211X1TF U461 ( .A0(N222), .A1(OPER_B[10]), .B0(N927), .C0(N928), .Y(N220)
         );
  AOI21X1TF U462 ( .A0(N975), .A1(N972), .B0(N910), .Y(N928) );
  AOI21X1TF U463 ( .A0(N926), .A1(N925), .B0(N924), .Y(N927) );
  AOI32X1TF U464 ( .A0(N923), .A1(OPER_B[10]), .A2(N922), .B0(N921), .B1(
        OPER_B[10]), .Y(N925) );
  AOI211X1TF U465 ( .A0(N920), .A1(OPER_B[11]), .B0(N919), .C0(N918), .Y(N926)
         );
  AOI21X1TF U466 ( .A0(N913), .A1(N917), .B0(N912), .Y(N914) );
  NOR3X1TF U467 ( .A(N911), .B(OPER_B[10]), .C(N923), .Y(N919) );
  AOI22X1TF U468 ( .A0(SUM_AB[4]), .A1(N87), .B0(N986), .B1(N1015), .Y(N987)
         );
  AOI22X1TF U469 ( .A0(DIVISION_HEAD[4]), .A1(N108), .B0(ZTEMP[4]), .B1(N141), 
        .Y(N988) );
  AOI22X1TF U470 ( .A0(SUM_AB[6]), .A1(N87), .B0(N992), .B1(N1015), .Y(N993)
         );
  AOI22X1TF U471 ( .A0(DIVISION_HEAD[6]), .A1(N108), .B0(ZTEMP[6]), .B1(N141), 
        .Y(N994) );
  AOI22X1TF U472 ( .A0(SUM_AB[2]), .A1(N87), .B0(N980), .B1(N1015), .Y(N981)
         );
  AOI22X1TF U473 ( .A0(DIVISION_HEAD[2]), .A1(N108), .B0(ZTEMP[2]), .B1(N141), 
        .Y(N982) );
  AOI22X1TF U474 ( .A0(SUM_AB[8]), .A1(N87), .B0(N998), .B1(N1015), .Y(N999)
         );
  AOI22X1TF U475 ( .A0(DIVISION_HEAD[8]), .A1(N108), .B0(ZTEMP[8]), .B1(N141), 
        .Y(N1000) );
  AOI22X1TF U476 ( .A0(SUM_AB[1]), .A1(N87), .B0(N977), .B1(N1015), .Y(N978)
         );
  AOI22X1TF U477 ( .A0(DIVISION_HEAD[1]), .A1(N108), .B0(ZTEMP[1]), .B1(N141), 
        .Y(N979) );
  AOI211X1TF U478 ( .A0(OPER_B[6]), .A1(N885), .B0(N884), .C0(N883), .Y(N886)
         );
  AOI21X1TF U479 ( .A0(N913), .A1(N882), .B0(N912), .Y(N880) );
  OAI31X1TF U480 ( .A0(N911), .A1(OPER_B[6]), .A2(N879), .B0(N878), .Y(N884)
         );
  AOI21X1TF U481 ( .A0(OPER_B[7]), .A1(N877), .B0(N876), .Y(N878) );
  OAI21X1TF U482 ( .A0(N911), .A1(N875), .B0(N874), .Y(N885) );
  OAI22X1TF U483 ( .A0(N513), .A1(N485), .B0(N484), .B1(N529), .Y(N710) );
  AOI211X1TF U484 ( .A0(SUM_AB[9]), .A1(N135), .B0(N482), .C0(N481), .Y(N485)
         );
  OAI211X1TF U485 ( .A0(N1003), .A1(N507), .B0(N480), .C0(N479), .Y(N481) );
  OAI22X1TF U486 ( .A0(N178), .A1(N100), .B0(N488), .B1(N609), .Y(N482) );
  OAI22X1TF U487 ( .A0(N475), .A1(N474), .B0(N473), .B1(N178), .Y(N711) );
  AOI211X1TF U488 ( .A0(N998), .A1(N493), .B0(N470), .C0(N469), .Y(N474) );
  OAI211X1TF U489 ( .A0(N468), .A1(N609), .B0(N467), .C0(N466), .Y(N469) );
  AOI22X1TF U490 ( .A0(XTEMP[9]), .A1(N96), .B0(N800), .B1(SUM_AB[12]), .Y(
        N466) );
  NOR2X1TF U491 ( .A(DIVISION_HEAD[12]), .B(N472), .Y(N465) );
  AOI22X1TF U492 ( .A0(X_IN[8]), .A1(N464), .B0(INTADD_0_N1), .B1(N488), .Y(
        N472) );
  OAI22X1TF U493 ( .A0(N154), .A1(N100), .B0(N463), .B1(N98), .Y(N470) );
  AOI22X1TF U494 ( .A0(SUM_AB[10]), .A1(N88), .B0(N1004), .B1(N1015), .Y(N1005) );
  AOI22X1TF U495 ( .A0(DIVISION_HEAD[10]), .A1(N108), .B0(ZTEMP[10]), .B1(N141), .Y(N1006) );
  AOI32X1TF U496 ( .A0(N431), .A1(N460), .A2(N430), .B0(N475), .B1(N157), .Y(
        N715) );
  AOI211X1TF U497 ( .A0(N493), .A1(N986), .B0(N429), .C0(N428), .Y(N430) );
  AOI22X1TF U498 ( .A0(DIVISION_HEAD[9]), .A1(N95), .B0(N82), .B1(N102), .Y(
        N426) );
  OAI22X1TF U499 ( .A0(N423), .A1(N100), .B0(N157), .B1(N454), .Y(N429) );
  AOI32X1TF U500 ( .A0(N411), .A1(N460), .A2(N410), .B0(N475), .B1(N155), .Y(
        N717) );
  AOI211X1TF U501 ( .A0(DIVISION_HEAD[7]), .A1(N96), .B0(N409), .C0(N408), .Y(
        N410) );
  OAI211X1TF U502 ( .A0(N98), .A1(N750), .B0(N407), .C0(N406), .Y(N408) );
  AOI21X1TF U503 ( .A0(N493), .A1(N980), .B0(N405), .Y(N406) );
  AOI22X1TF U504 ( .A0(X_IN[1]), .A1(N444), .B0(N800), .B1(SUM_AB[6]), .Y(N407) );
  OAI21X1TF U505 ( .A0(N500), .A1(N749), .B0(N402), .Y(N409) );
  AOI22X1TF U506 ( .A0(X_IN[8]), .A1(N137), .B0(X_IN[7]), .B1(N102), .Y(N402)
         );
  AOI32X1TF U507 ( .A0(N392), .A1(N391), .A2(N390), .B0(N475), .B1(N391), .Y(
        N719) );
  OAI211X1TF U508 ( .A0(N388), .A1(N559), .B0(N387), .C0(N386), .Y(N389) );
  AOI22X1TF U509 ( .A0(X_IN[6]), .A1(N137), .B0(N106), .B1(N102), .Y(N386) );
  AOI22X1TF U510 ( .A0(DIVISION_HEAD[3]), .A1(N736), .B0(SUM_AB[0]), .B1(N380), 
        .Y(N392) );
  AOI32X1TF U511 ( .A0(N461), .A1(N460), .A2(N459), .B0(N475), .B1(N154), .Y(
        N712) );
  OAI211X1TF U512 ( .A0(N507), .A1(N997), .B0(N456), .C0(N455), .Y(N457) );
  AOI22X1TF U513 ( .A0(DIVISION_HEAD[12]), .A1(N95), .B0(X_IN[12]), .B1(N102), 
        .Y(N455) );
  AOI22X1TF U514 ( .A0(DIVISION_HEAD[11]), .A1(N806), .B0(DIVISION_HEAD[10]), 
        .B1(N131), .Y(N456) );
  OAI22X1TF U515 ( .A0(N463), .A1(N609), .B0(N559), .B1(N498), .Y(N458) );
  AOI32X1TF U516 ( .A0(N401), .A1(N460), .A2(N400), .B0(N475), .B1(N514), .Y(
        N718) );
  AOI211X1TF U517 ( .A0(N493), .A1(N977), .B0(N399), .C0(N398), .Y(N400) );
  OAI211X1TF U518 ( .A0(N559), .A1(N432), .B0(N397), .C0(N396), .Y(N398) );
  AOI21X1TF U519 ( .A0(DIVISION_HEAD[4]), .A1(N736), .B0(N395), .Y(N396) );
  OAI22X1TF U520 ( .A0(N514), .A1(N454), .B0(N750), .B1(N609), .Y(N395) );
  AOI22X1TF U521 ( .A0(DIVISION_HEAD[6]), .A1(N96), .B0(X_IN[7]), .B1(N137), 
        .Y(N397) );
  OAI22X1TF U522 ( .A0(N463), .A1(N394), .B0(N488), .B1(N749), .Y(N399) );
  AOI32X1TF U523 ( .A0(N799), .A1(N816), .A2(N798), .B0(N814), .B1(N174), .Y(
        N684) );
  AOI21X1TF U524 ( .A0(N797), .A1(N1004), .B0(N796), .Y(N798) );
  AOI22X1TF U525 ( .A0(DIVISION_HEAD[0]), .A1(N131), .B0(DIVISION_HEAD[1]), 
        .B1(N806), .Y(N793) );
  AOI22X1TF U526 ( .A0(Y_IN[10]), .A1(N791), .B0(N94), .B1(N137), .Y(N794) );
  AOI22X1TF U527 ( .A0(N800), .A1(SUM_AB[1]), .B0(SUM_AB[10]), .B1(N146), .Y(
        N799) );
  OAI22X1TF U528 ( .A0(N513), .A1(N496), .B0(N495), .B1(N161), .Y(N709) );
  AOI21X1TF U529 ( .A0(N493), .A1(N1004), .B0(N492), .Y(N496) );
  OAI211X1TF U530 ( .A0(N500), .A1(N609), .B0(N491), .C0(N490), .Y(N492) );
  AOI22X1TF U531 ( .A0(XTEMP[11]), .A1(N96), .B0(SUM_AB[10]), .B1(N134), .Y(
        N491) );
  AOI21X1TF U532 ( .A0(SUM_AB[10]), .A1(N486), .B0(N499), .Y(N1004) );
  AOI22X1TF U533 ( .A0(N196), .A1(N149), .B0(N781), .B1(N780), .Y(N686) );
  AOI211X1TF U534 ( .A0(DIVISION_REMA[7]), .A1(N736), .B0(N779), .C0(N778), 
        .Y(N781) );
  OAI211X1TF U535 ( .A0(N173), .A1(N777), .B0(N776), .C0(N775), .Y(N778) );
  AOI22X1TF U536 ( .A0(N774), .A1(N773), .B0(N998), .B1(N797), .Y(N775) );
  AOI21X1TF U537 ( .A0(SUM_AB[8]), .A1(N462), .B0(N477), .Y(N998) );
  AOI32X1TF U538 ( .A0(N772), .A1(N771), .A2(N770), .B0(N769), .B1(N771), .Y(
        N773) );
  AOI22X1TF U539 ( .A0(DIVISION_REMA[8]), .A1(N763), .B0(SUM_AB[8]), .B1(N145), 
        .Y(N776) );
  AOI22X1TF U540 ( .A0(N475), .A1(N158), .B0(N441), .B1(N460), .Y(N714) );
  AOI21X1TF U541 ( .A0(DIVISION_HEAD[8]), .A1(N131), .B0(N434), .Y(N435) );
  OAI22X1TF U542 ( .A0(N158), .A1(N454), .B0(N507), .B1(N991), .Y(N434) );
  AOI22X1TF U543 ( .A0(DIVISION_HEAD[10]), .A1(N95), .B0(X_IN[10]), .B1(N101), 
        .Y(N437) );
  OAI22X1TF U544 ( .A0(N442), .A1(N609), .B0(N559), .B1(N476), .Y(N440) );
  AOI32X1TF U545 ( .A0(N421), .A1(N460), .A2(N420), .B0(N475), .B1(N423), .Y(
        N716) );
  AOI211X1TF U546 ( .A0(DIVISION_HEAD[8]), .A1(N96), .B0(N419), .C0(N418), .Y(
        N420) );
  OAI211X1TF U547 ( .A0(N559), .A1(N452), .B0(N417), .C0(N416), .Y(N418) );
  AOI21X1TF U548 ( .A0(DIVISION_HEAD[6]), .A1(N736), .B0(N415), .Y(N416) );
  OAI22X1TF U549 ( .A0(N423), .A1(N454), .B0(N507), .B1(N985), .Y(N415) );
  OAI21X1TF U550 ( .A0(N502), .A1(N749), .B0(N412), .Y(N419) );
  AOI22X1TF U551 ( .A0(X_IN[8]), .A1(N102), .B0(N82), .B1(N137), .Y(N412) );
  OAI211X1TF U552 ( .A0(N1010), .A1(N1009), .B0(N1008), .C0(N1007), .Y(N658)
         );
  AOI22X1TF U553 ( .A0(DIVISION_HEAD[11]), .A1(N108), .B0(ZTEMP[11]), .B1(N141), .Y(N1008) );
  OAI211X1TF U554 ( .A0(N1019), .A1(N1018), .B0(N1017), .C0(N1016), .Y(N657)
         );
  AOI32X1TF U555 ( .A0(N1018), .A1(N1015), .A2(N1014), .B0(N1013), .B1(N1015), 
        .Y(N1016) );
  AOI211X4TF U556 ( .A0(N975), .A1(N974), .B0(N973), .C0(N1011), .Y(N1015) );
  INVX2TF U557 ( .A(N970), .Y(N973) );
  AOI22X1TF U558 ( .A0(DIVISION_HEAD[12]), .A1(N108), .B0(ZTEMP[12]), .B1(
        N1011), .Y(N1017) );
  OAI31X1TF U559 ( .A0(N967), .A1(N61), .A2(N972), .B0(N966), .Y(N968) );
  AOI31X1TF U560 ( .A0(N182), .A1(N61), .A2(N965), .B0(N964), .Y(N966) );
  INVX2TF U561 ( .A(N1011), .Y(N969) );
  AOI31X1TF U562 ( .A0(N960), .A1(N959), .A2(N958), .B0(N957), .Y(N963) );
  OAI31X1TF U563 ( .A0(N956), .A1(N955), .A2(N954), .B0(N953), .Y(N957) );
  INVX2TF U564 ( .A(N922), .Y(N911) );
  OAI22X1TF U565 ( .A0(N513), .A1(N512), .B0(N511), .B1(N159), .Y(N708) );
  OAI21X1TF U566 ( .A0(N507), .A1(N1009), .B0(N506), .Y(N508) );
  AOI211X1TF U567 ( .A0(SUM_AB[11]), .A1(N134), .B0(N504), .C0(N503), .Y(N506)
         );
  INVX2TF U568 ( .A(N493), .Y(N507) );
  OAI21X1TF U569 ( .A0(N761), .A1(N183), .B0(N563), .Y(N705) );
  OAI22X1TF U570 ( .A0(N562), .A1(N561), .B0(N763), .B1(N780), .Y(N563) );
  AOI22X1TF U571 ( .A0(Y_IN[0]), .A1(N791), .B0(DIVISION_REMA[1]), .B1(N120), 
        .Y(N560) );
  AOI21X1TF U572 ( .A0(N119), .A1(N651), .B0(N976), .Y(N562) );
  INVX2TF U573 ( .A(SUM_AB[0]), .Y(N976) );
  OAI22X1TF U574 ( .A0(N196), .A1(N655), .B0(N761), .B1(N184), .Y(N693) );
  AOI21X1TF U575 ( .A0(SUM_AB[1]), .A1(N146), .B0(N654), .Y(N655) );
  AOI22X1TF U576 ( .A0(DIVISION_REMA[0]), .A1(N736), .B0(N797), .B1(N977), .Y(
        N652) );
  AOI21X1TF U577 ( .A0(SUM_AB[1]), .A1(SUM_AB[0]), .B0(N403), .Y(N977) );
  AOI22X1TF U578 ( .A0(Y_IN[1]), .A1(N791), .B0(DIVISION_REMA[2]), .B1(N125), 
        .Y(N653) );
  OAI22X1TF U579 ( .A0(N196), .A1(N741), .B0(N761), .B1(N175), .Y(N690) );
  AOI211X1TF U580 ( .A0(SUM_AB[4]), .A1(N146), .B0(N740), .C0(N739), .Y(N741)
         );
  OAI211X1TF U581 ( .A0(N738), .A1(N98), .B0(N757), .C0(N737), .Y(N739) );
  AOI22X1TF U582 ( .A0(DIVISION_REMA[5]), .A1(N125), .B0(N797), .B1(N986), .Y(
        N737) );
  AOI21X1TF U583 ( .A0(SUM_AB[4]), .A1(N422), .B0(N433), .Y(N986) );
  OAI22X1TF U584 ( .A0(N206), .A1(N804), .B0(N170), .B1(N100), .Y(N740) );
  OAI22X1TF U585 ( .A0(N196), .A1(N730), .B0(N761), .B1(N150), .Y(N692) );
  AOI211X1TF U586 ( .A0(SUM_AB[2]), .A1(N146), .B0(N729), .C0(N728), .Y(N730)
         );
  OAI211X1TF U587 ( .A0(N727), .A1(N98), .B0(N757), .C0(N656), .Y(N728) );
  AOI22X1TF U588 ( .A0(DIVISION_REMA[3]), .A1(N125), .B0(N797), .B1(N980), .Y(
        N656) );
  AOI21X1TF U589 ( .A0(SUM_AB[2]), .A1(N404), .B0(N414), .Y(N980) );
  NOR2X1TF U590 ( .A(SUM_AB[0]), .B(SUM_AB[1]), .Y(N403) );
  OAI22X1TF U591 ( .A0(N738), .A1(N804), .B0(N184), .B1(N100), .Y(N729) );
  OAI22X1TF U592 ( .A0(N196), .A1(N753), .B0(N761), .B1(N176), .Y(N688) );
  AOI211X1TF U593 ( .A0(N992), .A1(N797), .B0(N752), .C0(N751), .Y(N753) );
  OAI211X1TF U594 ( .A0(N750), .A1(N749), .B0(N757), .C0(N748), .Y(N751) );
  AOI22X1TF U595 ( .A0(DIVISION_REMA[7]), .A1(N120), .B0(SUM_AB[6]), .B1(N145), 
        .Y(N748) );
  INVX2TF U596 ( .A(N807), .Y(N749) );
  OAI21X1TF U597 ( .A0(N206), .A1(N98), .B0(N746), .Y(N752) );
  AOI22X1TF U598 ( .A0(Y_IN[6]), .A1(N791), .B0(DIVISION_REMA[5]), .B1(N736), 
        .Y(N746) );
  AOI21X1TF U599 ( .A0(SUM_AB[6]), .A1(N443), .B0(N453), .Y(N992) );
  OAI21X1TF U600 ( .A0(N761), .A1(N172), .B0(N760), .Y(N687) );
  OAI21X1TF U601 ( .A0(N759), .A1(N758), .B0(N780), .Y(N760) );
  INVX2TF U602 ( .A(N196), .Y(N780) );
  OAI211X1TF U603 ( .A0(N149), .A1(N777), .B0(N757), .C0(N756), .Y(N758) );
  AOI22X1TF U604 ( .A0(DIVISION_REMA[6]), .A1(N736), .B0(SUM_AB[7]), .B1(N145), 
        .Y(N756) );
  OAI211X1TF U605 ( .A0(N810), .A1(N997), .B0(N755), .C0(N754), .Y(N759) );
  OAI21X1TF U606 ( .A0(N453), .A1(N452), .B0(N462), .Y(N997) );
  OAI22X1TF U607 ( .A0(N513), .A1(N362), .B0(N361), .B1(N179), .Y(N723) );
  AOI211X1TF U608 ( .A0(N493), .A1(N1013), .B0(N359), .C0(N358), .Y(N362) );
  OAI31X1TF U609 ( .A0(XTEMP[12]), .A1(N360), .A2(N509), .B0(N357), .Y(N358)
         );
  AOI22X1TF U610 ( .A0(XTEMP[11]), .A1(N131), .B0(N139), .B1(N444), .Y(N357)
         );
  INVX2TF U611 ( .A(N609), .Y(N444) );
  NAND2X2TF U612 ( .A(MODE_TYPE[1]), .B(N356), .Y(N609) );
  INVX2TF U613 ( .A(INTADD_0_N1), .Y(N464) );
  NOR2X1TF U614 ( .A(N156), .B(N750), .Y(INTADD_0_CI) );
  INVX2TF U615 ( .A(X_IN[0]), .Y(N750) );
  OAI22X1TF U616 ( .A0(N119), .A1(N1018), .B0(N502), .B1(N98), .Y(N359) );
  NOR2X2TF U617 ( .A(N393), .B(N1018), .Y(N493) );
  AOI31X1TF U618 ( .A0(N941), .A1(N73), .A2(N564), .B0(N353), .Y(N384) );
  OAI211X1TF U619 ( .A0(N73), .A1(N378), .B0(N363), .C0(N352), .Y(N353) );
  OAI211X1TF U620 ( .A0(N960), .A1(N351), .B0(N567), .C0(N601), .Y(N352) );
  NOR2X1TF U621 ( .A(PRE_WORK), .B(N368), .Y(N603) );
  INVX2TF U622 ( .A(N600), .Y(N567) );
  NOR2X1TF U623 ( .A(N375), .B(N944), .Y(N363) );
  INVX2TF U624 ( .A(N393), .Y(N375) );
  INVX2TF U625 ( .A(N618), .Y(N378) );
  OAI22X1TF U626 ( .A0(N196), .A1(N735), .B0(N761), .B1(N170), .Y(N691) );
  AOI211X1TF U627 ( .A0(SUM_AB[3]), .A1(N146), .B0(N734), .C0(N733), .Y(N735)
         );
  OAI211X1TF U628 ( .A0(N810), .A1(N985), .B0(N757), .C0(N732), .Y(N733) );
  OAI21X1TF U629 ( .A0(N414), .A1(N413), .B0(N422), .Y(N985) );
  OAI22X1TF U630 ( .A0(N731), .A1(N804), .B0(N150), .B1(N100), .Y(N734) );
  OAI22X1TF U631 ( .A0(N196), .A1(N745), .B0(N761), .B1(N171), .Y(N689) );
  AOI211X1TF U632 ( .A0(SUM_AB[5]), .A1(N146), .B0(N744), .C0(N743), .Y(N745)
         );
  OAI211X1TF U633 ( .A0(N810), .A1(N991), .B0(N757), .C0(N742), .Y(N743) );
  AOI222X4TF U634 ( .A0(N767), .A1(N101), .B0(N765), .B1(N136), .C0(N558), 
        .C1(N807), .Y(N757) );
  OAI21X1TF U635 ( .A0(N433), .A1(N432), .B0(N443), .Y(N991) );
  INVX2TF U636 ( .A(N804), .Y(N791) );
  NOR3X1TF U637 ( .A(N774), .B(N131), .C(N557), .Y(N782) );
  AOI32X1TF U638 ( .A0(N790), .A1(N816), .A2(N789), .B0(N814), .B1(N173), .Y(
        N685) );
  OAI211X1TF U639 ( .A0(N810), .A1(N1003), .B0(N786), .C0(N785), .Y(N787) );
  AOI22X1TF U640 ( .A0(DIVISION_HEAD[1]), .A1(N125), .B0(X_IN[1]), .B1(N101), 
        .Y(N785) );
  OAI21X1TF U641 ( .A0(N477), .A1(N476), .B0(N486), .Y(N1003) );
  OAI21X1TF U642 ( .A0(N784), .A1(N804), .B0(N783), .Y(N788) );
  AOI22X1TF U643 ( .A0(DIVISION_REMA[8]), .A1(N131), .B0(N800), .B1(SUM_AB[0]), 
        .Y(N783) );
  AOI22X1TF U644 ( .A0(DIVISION_HEAD[0]), .A1(N806), .B0(SUM_AB[9]), .B1(N146), 
        .Y(N790) );
  AOI32X1TF U645 ( .A0(N817), .A1(N816), .A2(N815), .B0(N814), .B1(N167), .Y(
        N683) );
  AOI211X1TF U646 ( .A0(DIVISION_HEAD[3]), .A1(N125), .B0(N812), .C0(N811), 
        .Y(N815) );
  OAI211X1TF U647 ( .A0(N810), .A1(N1009), .B0(N809), .C0(N808), .Y(N811) );
  AOI22X1TF U648 ( .A0(DIVISION_HEAD[1]), .A1(N131), .B0(DIVISION_HEAD[2]), 
        .B1(N806), .Y(N809) );
  OAI21X1TF U649 ( .A0(N499), .A1(N498), .B0(N1014), .Y(N1009) );
  INVX2TF U650 ( .A(N797), .Y(N810) );
  OAI21X1TF U651 ( .A0(N805), .A1(N804), .B0(N803), .Y(N812) );
  INVX2TF U652 ( .A(N97), .Y(N802) );
  INVX2TF U653 ( .A(N814), .Y(N816) );
  AOI22X1TF U654 ( .A0(N800), .A1(SUM_AB[2]), .B0(SUM_AB[11]), .B1(N146), .Y(
        N817) );
  OAI21X1TF U655 ( .A0(N814), .A1(N556), .B0(N555), .Y(N706) );
  OAI21X1TF U656 ( .A0(N814), .A1(N806), .B0(DIVISION_HEAD[3]), .Y(N555) );
  INVX2TF U657 ( .A(N454), .Y(N806) );
  AOI211X1TF U658 ( .A0(DIVISION_HEAD[2]), .A1(N131), .B0(N554), .C0(N553), 
        .Y(N556) );
  AOI22X1TF U659 ( .A0(N800), .A1(SUM_AB[3]), .B0(N1013), .B1(N797), .Y(N550)
         );
  NOR2X2TF U660 ( .A(N1018), .B(N651), .Y(N797) );
  NOR2X1TF U661 ( .A(N1018), .B(N1014), .Y(N1013) );
  INVX2TF U662 ( .A(SUM_AB[11]), .Y(N498) );
  INVX2TF U663 ( .A(SUM_AB[9]), .Y(N476) );
  INVX2TF U664 ( .A(SUM_AB[7]), .Y(N452) );
  NOR2X1TF U665 ( .A(SUM_AB[6]), .B(N443), .Y(N453) );
  INVX2TF U666 ( .A(SUM_AB[5]), .Y(N432) );
  NOR2X1TF U667 ( .A(SUM_AB[4]), .B(N422), .Y(N433) );
  INVX2TF U668 ( .A(SUM_AB[3]), .Y(N413) );
  NOR3X1TF U669 ( .A(SUM_AB[0]), .B(SUM_AB[2]), .C(SUM_AB[1]), .Y(N414) );
  INVX2TF U670 ( .A(SUM_AB[12]), .Y(N1018) );
  INVX2TF U671 ( .A(N559), .Y(N800) );
  AOI22X1TF U672 ( .A0(N941), .A1(SUM_AB[12]), .B0(N106), .B1(N137), .Y(N551)
         );
  OAI21X1TF U673 ( .A0(N179), .A1(N112), .B0(N260), .Y(OPER_A[12]) );
  AND2X2TF U674 ( .A(N764), .B(N769), .Y(N766) );
  INVX2TF U675 ( .A(N385), .Y(N774) );
  OAI22X1TF U676 ( .A0(N549), .A1(N804), .B0(N548), .B1(N98), .Y(N554) );
  NAND2X2TF U677 ( .A(N356), .B(N315), .Y(N804) );
  INVX2TF U678 ( .A(N356), .Y(N640) );
  AOI31X1TF U679 ( .A0(N122), .A1(N383), .A2(N382), .B0(N381), .Y(N547) );
  INVX2TF U680 ( .A(N308), .Y(N765) );
  OAI211X1TF U681 ( .A0(X_IN[12]), .A1(N548), .B0(N307), .C0(N306), .Y(N308)
         );
  OAI22X1TF U682 ( .A0(Y_IN[10]), .A1(N305), .B0(N304), .B1(N303), .Y(N306) );
  OAI22X1TF U683 ( .A0(X_IN[10]), .A1(N302), .B0(N138), .B1(N784), .Y(N303) );
  OAI21X1TF U684 ( .A0(Y_IN[9]), .A1(N201), .B0(Y_IN[8]), .Y(N302) );
  AOI211X1TF U685 ( .A0(X_IN[10]), .A1(N762), .B0(N301), .C0(N300), .Y(N304)
         );
  AOI21X1TF U686 ( .A0(N89), .A1(N500), .B0(N299), .Y(N300) );
  AOI211X1TF U687 ( .A0(X_IN[8]), .A1(N298), .B0(N297), .C0(N296), .Y(N299) );
  NOR2X1TF U688 ( .A(N89), .B(N500), .Y(N297) );
  AOI21X1TF U689 ( .A0(N197), .A1(N468), .B0(N295), .Y(N298) );
  AOI211X1TF U690 ( .A0(X_IN[6]), .A1(N294), .B0(N293), .C0(N292), .Y(N295) );
  NOR2X1TF U691 ( .A(N197), .B(N468), .Y(N293) );
  AOI32X1TF U692 ( .A0(N291), .A1(N290), .A2(N319), .B0(N289), .B1(N290), .Y(
        N294) );
  OAI22X1TF U693 ( .A0(X_IN[4]), .A1(N738), .B0(N106), .B1(N731), .Y(N289) );
  OAI32X1TF U694 ( .A0(N288), .A1(N93), .A2(N317), .B0(X_IN[2]), .B1(N288), 
        .Y(N291) );
  INVX2TF U695 ( .A(X_IN[7]), .Y(N468) );
  INVX2TF U696 ( .A(X_IN[9]), .Y(N500) );
  NOR2X1TF U697 ( .A(Y_IN[9]), .B(N201), .Y(N301) );
  NOR2X1TF U698 ( .A(Y_IN[12]), .B(Y_IN[11]), .Y(N307) );
  INVX2TF U699 ( .A(N770), .Y(N558) );
  OR2X2TF U700 ( .A(MODE_TYPE[0]), .B(N315), .Y(N769) );
  INVX2TF U701 ( .A(MODE_TYPE[1]), .Y(N315) );
  OAI31X1TF U702 ( .A0(N286), .A1(N139), .A2(N548), .B0(N285), .Y(N287) );
  OAI31X1TF U703 ( .A0(N284), .A1(N283), .A2(N282), .B0(N281), .Y(N285) );
  AOI22X1TF U704 ( .A0(N138), .A1(N548), .B0(X_IN[12]), .B1(N805), .Y(N281) );
  NOR2X1TF U705 ( .A(X_IN[10]), .B(N784), .Y(N282) );
  AOI211X1TF U706 ( .A0(X_IN[10]), .A1(N784), .B0(X_IN[9]), .C0(N762), .Y(N283) );
  AOI211X1TF U707 ( .A0(X_IN[9]), .A1(N762), .B0(N280), .C0(N279), .Y(N284) );
  AOI21X1TF U708 ( .A0(N89), .A1(N488), .B0(N278), .Y(N279) );
  AOI211X1TF U709 ( .A0(N277), .A1(X_IN[7]), .B0(N276), .C0(N275), .Y(N278) );
  NOR2X1TF U710 ( .A(N89), .B(N488), .Y(N276) );
  AOI21X1TF U711 ( .A0(N197), .A1(N463), .B0(N274), .Y(N277) );
  AOI211X1TF U712 ( .A0(N273), .A1(N106), .B0(N272), .C0(N271), .Y(N274) );
  NOR2X1TF U713 ( .A(N197), .B(N463), .Y(N272) );
  AOI211X1TF U714 ( .A0(Y_IN[3]), .A1(N442), .B0(N270), .C0(N269), .Y(N273) );
  AOI211X1TF U715 ( .A0(X_IN[4]), .A1(N731), .B0(N94), .C0(N738), .Y(N269) );
  OAI32X1TF U716 ( .A0(N268), .A1(X_IN[2]), .A2(N317), .B0(X_IN[1]), .B1(N268), 
        .Y(N270) );
  OAI211X1TF U717 ( .A0(Y_IN[3]), .A1(N442), .B0(N267), .C0(N319), .Y(N268) );
  AOI22X1TF U718 ( .A0(N93), .A1(N738), .B0(X_IN[2]), .B1(N318), .Y(N267) );
  INVX2TF U719 ( .A(X_IN[4]), .Y(N442) );
  INVX2TF U720 ( .A(X_IN[6]), .Y(N463) );
  INVX2TF U721 ( .A(X_IN[8]), .Y(N488) );
  NOR2X1TF U722 ( .A(Y_IN[9]), .B(N502), .Y(N280) );
  INVX2TF U723 ( .A(X_IN[10]), .Y(N502) );
  NOR2X1TF U724 ( .A(Y_IN[11]), .B(N305), .Y(N286) );
  INVX2TF U725 ( .A(X_IN[12]), .Y(N305) );
  INVX2TF U726 ( .A(N342), .Y(N383) );
  OAI211X1TF U727 ( .A0(N862), .A1(N861), .B0(N860), .C0(N859), .Y(N678) );
  AOI32X1TF U728 ( .A0(N937), .A1(OPER_B[4]), .A2(N858), .B0(N890), .B1(
        OPER_B[4]), .Y(N859) );
  AOI211X1TF U729 ( .A0(N864), .A1(OPER_B[5]), .B0(N857), .C0(N856), .Y(N860)
         );
  OAI31X1TF U730 ( .A0(N934), .A1(OPER_A[4]), .A2(N855), .B0(N210), .Y(N856)
         );
  AOI21X1TF U731 ( .A0(N113), .A1(C152_DATA4_4), .B0(N211), .Y(N210) );
  NOR3X1TF U732 ( .A(OPER_B[4]), .B(N858), .C(N116), .Y(N857) );
  AOI21X1TF U733 ( .A0(N931), .A1(N855), .B0(N854), .Y(N861) );
  OAI211X1TF U734 ( .A0(N830), .A1(N832), .B0(N829), .C0(N212), .Y(N681) );
  AOI211X1TF U735 ( .A0(N114), .A1(C152_DATA4_1), .B0(N826), .C0(N891), .Y(
        N212) );
  OAI31X1TF U736 ( .A0(OPER_B[1]), .A1(N116), .A2(N189), .B0(N825), .Y(N826)
         );
  AOI211X1TF U737 ( .A0(N864), .A1(OPER_B[2]), .B0(N828), .C0(N827), .Y(N829)
         );
  NOR3X1TF U738 ( .A(N831), .B(OPER_A[1]), .C(N934), .Y(N827) );
  OAI32X1TF U739 ( .A0(N187), .A1(OPER_B[0]), .A2(N116), .B0(N935), .B1(N187), 
        .Y(N828) );
  AOI21X1TF U740 ( .A0(N931), .A1(N831), .B0(N854), .Y(N830) );
  INVX2TF U741 ( .A(N932), .Y(N854) );
  AOI211X1TF U742 ( .A0(N114), .A1(C152_DATA4_5), .B0(N866), .C0(N215), .Y(
        N216) );
  OAI31X1TF U743 ( .A0(OPER_B[5]), .A1(N865), .A2(N116), .B0(N905), .Y(N866)
         );
  OAI211X1TF U744 ( .A0(SIGN_Y), .A1(N965), .B0(N225), .C0(N972), .Y(N905) );
  AOI22X1TF U745 ( .A0(N864), .A1(OPER_B[6]), .B0(N863), .B1(N868), .Y(N873)
         );
  NOR2X1TF U746 ( .A(N934), .B(OPER_A[5]), .Y(N863) );
  INVX2TF U747 ( .A(N894), .Y(N864) );
  AOI22X1TF U748 ( .A0(OPER_B[5]), .A1(N870), .B0(OPER_A[5]), .B1(N869), .Y(
        N872) );
  OAI21X1TF U749 ( .A0(N934), .A1(N868), .B0(N932), .Y(N869) );
  OAI21X1TF U750 ( .A0(N116), .A1(N867), .B0(N935), .Y(N870) );
  OR2X2TF U751 ( .A(N930), .B(N891), .Y(N211) );
  NOR2X1TF U752 ( .A(N967), .B(N836), .Y(N876) );
  INVX2TF U753 ( .A(N935), .Y(N890) );
  NOR3X1TF U754 ( .A(N73), .B(N182), .C(N965), .Y(N964) );
  OAI22X1TF U755 ( .A0(N133), .A1(N206), .B0(OFFSET[2]), .B1(N207), .Y(C2_Z_4)
         );
  INVX2TF U756 ( .A(Y_IN[4]), .Y(N206) );
  OAI22X1TF U757 ( .A0(N133), .A1(N205), .B0(OFFSET[3]), .B1(N207), .Y(C2_Z_5)
         );
  OAI22X1TF U758 ( .A0(N132), .A1(N204), .B0(OFFSET[4]), .B1(N207), .Y(C2_Z_6)
         );
  OAI22X1TF U759 ( .A0(N132), .A1(N198), .B0(OFFSET[5]), .B1(N207), .Y(C2_Z_7)
         );
  INVX2TF U760 ( .A(Y_IN[11]), .Y(N805) );
  NOR2X1TF U761 ( .A(OPER_B[9]), .B(N908), .Y(N923) );
  NOR2X1TF U762 ( .A(N875), .B(OPER_B[6]), .Y(N892) );
  INVX2TF U763 ( .A(N879), .Y(N875) );
  NOR2X1TF U764 ( .A(OPER_B[5]), .B(N867), .Y(N879) );
  NOR2X1TF U765 ( .A(OPER_B[3]), .B(N847), .Y(N858) );
  AOI211X1TF U766 ( .A0(N61), .A1(N965), .B0(SIGN_Y), .C0(N910), .Y(N930) );
  NOR2X1TF U767 ( .A(OPER_A[9]), .B(N909), .Y(N917) );
  NOR2X1TF U768 ( .A(OPER_A[7]), .B(N893), .Y(N898) );
  NOR2X1TF U769 ( .A(OPER_A[5]), .B(N868), .Y(N882) );
  NOR2X1TF U770 ( .A(OPER_A[3]), .B(N846), .Y(N855) );
  OAI21X1TF U771 ( .A0(N157), .A1(N112), .B0(N251), .Y(OPER_A[4]) );
  OAI21X1TF U772 ( .A0(N158), .A1(N112), .B0(N252), .Y(OPER_A[5]) );
  OAI21X1TF U773 ( .A0(N160), .A1(N112), .B0(N253), .Y(OPER_A[6]) );
  OAI21X1TF U774 ( .A0(N154), .A1(N112), .B0(N254), .Y(OPER_A[7]) );
  OAI21X1TF U775 ( .A0(N178), .A1(N112), .B0(N255), .Y(OPER_A[8]) );
  OAI21X1TF U776 ( .A0(N112), .A1(N529), .B0(N256), .Y(OPER_A[9]) );
  OAI21X1TF U777 ( .A0(N112), .A1(N161), .B0(N257), .Y(OPER_A[10]) );
  OAI21X1TF U778 ( .A0(N112), .A1(N159), .B0(N258), .Y(OPER_A[11]) );
  OAI211X1TF U779 ( .A0(N181), .A1(N938), .B0(N853), .C0(N852), .Y(N679) );
  AOI211X1TF U780 ( .A0(OPER_A[3]), .A1(N851), .B0(N850), .C0(N849), .Y(N852)
         );
  OAI31X1TF U781 ( .A0(N934), .A1(OPER_A[3]), .A2(N848), .B0(N209), .Y(N849)
         );
  AOI21X1TF U782 ( .A0(C152_DATA4_3), .A1(N113), .B0(N906), .Y(N209) );
  NOR2X1TF U783 ( .A(N61), .B(N910), .Y(N906) );
  OAI21X1TF U784 ( .A0(N133), .A1(N317), .B0(N207), .Y(C2_Z_1) );
  OAI22X1TF U785 ( .A0(N133), .A1(N731), .B0(OFFSET[1]), .B1(N207), .Y(C2_Z_3)
         );
  INVX2TF U786 ( .A(Y_IN[3]), .Y(N731) );
  OAI32X1TF U787 ( .A0(N188), .A1(N115), .A2(N847), .B0(N935), .B1(N188), .Y(
        N850) );
  INVX2TF U788 ( .A(N874), .Y(N921) );
  AOI32X1TF U789 ( .A0(N606), .A1(N350), .A2(N824), .B0(N946), .B1(N349), .Y(
        N874) );
  INVX2TF U790 ( .A(N940), .Y(N946) );
  OAI21X1TF U791 ( .A0(N934), .A1(N846), .B0(N932), .Y(N851) );
  INVX2TF U792 ( .A(N837), .Y(N912) );
  AOI21X1TF U793 ( .A0(N565), .A1(N349), .B0(N564), .Y(N837) );
  INVX2TF U794 ( .A(N848), .Y(N846) );
  NOR3X1TF U795 ( .A(OPER_A[2]), .B(OPER_A[1]), .C(OPER_A[0]), .Y(N848) );
  OAI21X1TF U796 ( .A0(N155), .A1(N111), .B0(N249), .Y(OPER_A[2]) );
  INVX2TF U797 ( .A(N931), .Y(N934) );
  NOR2X2TF U798 ( .A(N924), .B(N916), .Y(N931) );
  INVX2TF U799 ( .A(N904), .Y(N924) );
  OAI21X1TF U800 ( .A0(N423), .A1(N111), .B0(N250), .Y(OPER_A[3]) );
  AOI31X1TF U801 ( .A0(N937), .A1(N188), .A2(N847), .B0(N888), .Y(N853) );
  OAI21X1TF U802 ( .A0(N975), .A1(N910), .B0(N843), .Y(N888) );
  INVX2TF U803 ( .A(N910), .Y(N225) );
  INVX2TF U804 ( .A(N348), .Y(N959) );
  INVX2TF U805 ( .A(N566), .Y(N949) );
  NOR2X1TF U806 ( .A(OPER_B[1]), .B(OPER_B[0]), .Y(N839) );
  INVX2TF U807 ( .A(N349), .Y(N350) );
  INVX2TF U808 ( .A(N606), .Y(N823) );
  NOR2X2TF U809 ( .A(N604), .B(N632), .Y(N824) );
  AOI221X1TF U810 ( .A0(N128), .A1(N164), .B0(N186), .B1(N91), .C0(N819), .Y(
        N820) );
  AOI22X1TF U811 ( .A0(\INDEX[2] ), .A1(N90), .B0(N124), .B1(\RSHT_BITS[3] ), 
        .Y(N818) );
  AOI32X1TF U812 ( .A0(N940), .A1(N953), .A2(N372), .B0(N955), .B1(N953), .Y(
        N346) );
  OR2X2TF U813 ( .A(N632), .B(N152), .Y(N372) );
  INVX2TF U814 ( .A(N604), .Y(N643) );
  OAI21X1TF U815 ( .A0(N348), .A1(N939), .B0(N344), .Y(N608) );
  OAI21X1TF U816 ( .A0(N571), .A1(N565), .B0(N345), .Y(N344) );
  NOR2X2TF U817 ( .A(\RSHT_BITS[3] ), .B(N592), .Y(N606) );
  NOR3X1TF U818 ( .A(N121), .B(N122), .C(N954), .Y(N822) );
  INVX2TF U819 ( .A(N960), .Y(N967) );
  NOR2X1TF U820 ( .A(SIGN_Y), .B(N117), .Y(N907) );
  INVX2TF U821 ( .A(N312), .Y(N628) );
  OAI22X1TF U822 ( .A0(Y_IN[12]), .A1(N178), .B0(N340), .B1(N339), .Y(N341) );
  OAI31X1TF U823 ( .A0(N338), .A1(DIVISION_HEAD[10]), .A2(N548), .B0(N337), 
        .Y(N339) );
  AOI22X1TF U824 ( .A0(Y_IN[11]), .A1(N154), .B0(N336), .B1(N335), .Y(N337) );
  OAI22X1TF U825 ( .A0(DIVISION_HEAD[8]), .A1(N762), .B0(DIVISION_HEAD[9]), 
        .B1(N784), .Y(N335) );
  INVX2TF U826 ( .A(N334), .Y(N336) );
  NOR2X1TF U827 ( .A(Y_IN[11]), .B(N154), .Y(N338) );
  AOI211X1TF U828 ( .A0(DIVISION_HEAD[8]), .A1(N762), .B0(N333), .C0(N334), 
        .Y(N340) );
  OAI21X1TF U829 ( .A0(Y_IN[11]), .A1(N154), .B0(N332), .Y(N334) );
  AOI22X1TF U830 ( .A0(DIVISION_HEAD[10]), .A1(N548), .B0(DIVISION_HEAD[9]), 
        .B1(N784), .Y(N332) );
  INVX2TF U831 ( .A(Y_IN[9]), .Y(N784) );
  INVX2TF U832 ( .A(Y_IN[10]), .Y(N548) );
  AOI21X1TF U833 ( .A0(N89), .A1(N423), .B0(N331), .Y(N333) );
  AOI211X1TF U834 ( .A0(N330), .A1(DIVISION_HEAD[6]), .B0(N329), .C0(N328), 
        .Y(N331) );
  NOR2X1TF U835 ( .A(N89), .B(N423), .Y(N329) );
  AOI211X1TF U836 ( .A0(N326), .A1(DIVISION_HEAD[4]), .B0(N325), .C0(N324), 
        .Y(N327) );
  NOR2X1TF U837 ( .A(Y_IN[5]), .B(N514), .Y(N325) );
  AOI21X1TF U838 ( .A0(Y_IN[3]), .A1(N649), .B0(N323), .Y(N326) );
  OAI32X1TF U839 ( .A0(N322), .A1(DIVISION_HEAD[2]), .A2(N738), .B0(N321), 
        .B1(N322), .Y(N323) );
  OAI211X1TF U840 ( .A0(Y_IN[2]), .A1(N167), .B0(N320), .C0(N319), .Y(N321) );
  INVX2TF U841 ( .A(Y_IN[0]), .Y(N727) );
  INVX2TF U842 ( .A(Y_IN[1]), .Y(N317) );
  INVX2TF U843 ( .A(Y_IN[2]), .Y(N738) );
  INVX2TF U844 ( .A(Y_IN[8]), .Y(N762) );
  INVX2TF U845 ( .A(Y_IN[12]), .Y(N549) );
  NOR2X1TF U846 ( .A(N104), .B(N179), .Y(FOUT[12]) );
  NOR2X1TF U847 ( .A(N104), .B(N159), .Y(FOUT[11]) );
  OAI21X1TF U848 ( .A0(N178), .A1(N104), .B0(N243), .Y(FOUT[8]) );
  AOI21X1TF U849 ( .A0(N224), .A1(DIVISION_REMA[8]), .B0(N242), .Y(N243) );
  OAI22X1TF U850 ( .A0(N174), .A1(N86), .B0(N161), .B1(N84), .Y(N242) );
  OAI21X1TF U851 ( .A0(N154), .A1(N104), .B0(N241), .Y(FOUT[7]) );
  AOI21X1TF U852 ( .A0(N224), .A1(DIVISION_REMA[7]), .B0(N240), .Y(N241) );
  OAI22X1TF U853 ( .A0(N173), .A1(N86), .B0(N529), .B1(N84), .Y(N240) );
  OAI21X1TF U854 ( .A0(N160), .A1(N104), .B0(N239), .Y(FOUT[6]) );
  AOI21X1TF U855 ( .A0(N224), .A1(DIVISION_REMA[6]), .B0(N238), .Y(N239) );
  OAI22X1TF U856 ( .A0(N178), .A1(N84), .B0(N149), .B1(N86), .Y(N238) );
  OAI21X1TF U857 ( .A0(N514), .A1(N103), .B0(N229), .Y(FOUT[1]) );
  AOI21X1TF U858 ( .A0(N224), .A1(DIVISION_REMA[1]), .B0(N228), .Y(N229) );
  OAI22X1TF U859 ( .A0(N423), .A1(N83), .B0(N170), .B1(N85), .Y(N228) );
  OAI21X1TF U860 ( .A0(N158), .A1(N103), .B0(N237), .Y(FOUT[5]) );
  AOI21X1TF U861 ( .A0(N224), .A1(DIVISION_REMA[5]), .B0(N236), .Y(N237) );
  OAI22X1TF U862 ( .A0(N154), .A1(N83), .B0(N172), .B1(N85), .Y(N236) );
  OAI21X1TF U863 ( .A0(N155), .A1(N103), .B0(N231), .Y(FOUT[2]) );
  AOI21X1TF U864 ( .A0(N224), .A1(DIVISION_REMA[2]), .B0(N230), .Y(N231) );
  OAI22X1TF U865 ( .A0(N157), .A1(N83), .B0(N175), .B1(N85), .Y(N230) );
  OAI21X1TF U866 ( .A0(N157), .A1(N103), .B0(N235), .Y(FOUT[4]) );
  AOI21X1TF U867 ( .A0(N224), .A1(DIVISION_REMA[4]), .B0(N234), .Y(N235) );
  OAI22X1TF U868 ( .A0(N160), .A1(N83), .B0(N176), .B1(N85), .Y(N234) );
  OAI21X1TF U869 ( .A0(N423), .A1(N103), .B0(N233), .Y(FOUT[3]) );
  AOI21X1TF U870 ( .A0(N224), .A1(DIVISION_REMA[3]), .B0(N232), .Y(N233) );
  OAI22X1TF U871 ( .A0(N158), .A1(N83), .B0(N171), .B1(N85), .Y(N232) );
  NOR2X1TF U872 ( .A(N342), .B(N373), .Y(ALU_IS_DONE) );
  OAI211X1TF U873 ( .A0(N155), .A1(N84), .B0(N227), .C0(N226), .Y(FOUT[0]) );
  AOI22X1TF U874 ( .A0(N127), .A1(\INTADD_0_SUM[5] ), .B0(N800), .B1(
        SUM_AB[10]), .Y(N448) );
  AOI21X1TF U875 ( .A0(N127), .A1(N472), .B0(N471), .Y(N473) );
  AOI22X1TF U876 ( .A0(N126), .A1(N465), .B0(SUM_AB[8]), .B1(N134), .Y(N467)
         );
  AOI22X1TF U877 ( .A0(N127), .A1(\INTADD_0_SUM[3] ), .B0(SUM_AB[4]), .B1(N135), .Y(N431) );
  AOI22X1TF U878 ( .A0(N127), .A1(\INTADD_0_SUM[1] ), .B0(SUM_AB[2]), .B1(N135), .Y(N411) );
  AOI31X1TF U879 ( .A0(X_IN[0]), .A1(N127), .A2(N156), .B0(N389), .Y(N390) );
  AOI22X1TF U880 ( .A0(N127), .A1(\INTADD_0_SUM[6] ), .B0(SUM_AB[7]), .B1(N135), .Y(N461) );
  AOI22X1TF U881 ( .A0(N127), .A1(\INTADD_0_SUM[0] ), .B0(SUM_AB[1]), .B1(N135), .Y(N401) );
  AOI31X1TF U882 ( .A0(N126), .A1(N161), .A2(N494), .B0(N489), .Y(N490) );
  AOI22X1TF U883 ( .A0(N126), .A1(\INTADD_0_SUM[4] ), .B0(SUM_AB[5]), .B1(N134), .Y(N438) );
  AOI22X1TF U884 ( .A0(N127), .A1(\INTADD_0_SUM[2] ), .B0(SUM_AB[3]), .B1(N135), .Y(N421) );
  AOI31X1TF U885 ( .A0(N127), .A1(N159), .A2(N510), .B0(N508), .Y(N512) );
  AOI21X1TF U886 ( .A0(N127), .A1(N360), .B0(N513), .Y(N361) );
  NAND3X1TF U887 ( .A(N905), .B(N219), .C(N218), .Y(N674) );
  NAND4BX1TF U888 ( .AN(N844), .B(N214), .C(N845), .D(N213), .Y(N680) );
  AOI2BB2X1TF U889 ( .B0(N114), .B1(C152_DATA4_2), .A0N(N162), .A1N(N929), .Y(
        N213) );
  OAI2BB1X1TF U890 ( .A0N(N114), .A1N(C152_DATA4_10), .B0(N220), .Y(N672) );
  NAND3X1TF U891 ( .A(N872), .B(N873), .C(N216), .Y(N677) );
  OAI2BB2XLTF U892 ( .B0(OFFSET[0]), .B1(N207), .A0N(Y_IN[2]), .A1N(N81), .Y(
        C2_Z_2) );
  AOI2BB2X1TF U893 ( .B0(N224), .B1(DIVISION_REMA[0]), .A0N(N150), .A1N(N86), 
        .Y(N227) );
  OAI222X1TF U894 ( .A0(N84), .A1(N179), .B0(N86), .B1(N649), .C0(N104), .C1(
        N161), .Y(FOUT[10]) );
  OAI222X1TF U895 ( .A0(N104), .A1(N529), .B0(N86), .B1(N167), .C0(N159), .C1(
        N84), .Y(FOUT[9]) );
  NAND2X1TF U896 ( .A(N152), .B(N169), .Y(N373) );
  NAND3X1TF U897 ( .A(STEP[2]), .B(STEP[3]), .C(N643), .Y(N940) );
  NAND3X1TF U898 ( .A(N546), .B(N385), .C(N635), .Y(N648) );
  NOR4XLTF U899 ( .A(N763), .B(N618), .C(N802), .D(N648), .Y(N266) );
  AOI222XLTF U900 ( .A0(STEP[2]), .A1(N153), .B0(N121), .B1(N169), .C0(N151), 
        .C1(N122), .Y(N264) );
  NAND3X1TF U901 ( .A(N266), .B(N364), .C(N634), .Y(N620) );
  AOI2BB1X1TF U902 ( .A0N(N106), .A1N(N273), .B0(Y_IN[4]), .Y(N271) );
  AOI2BB1X1TF U903 ( .A0N(X_IN[7]), .A1N(N277), .B0(Y_IN[6]), .Y(N275) );
  NAND2X1TF U904 ( .A(MODE_TYPE[0]), .B(N315), .Y(N764) );
  AO22X1TF U905 ( .A0(X_IN[4]), .A1(N738), .B0(N93), .B1(N318), .Y(N288) );
  NAND2X1TF U906 ( .A(N105), .B(N731), .Y(N290) );
  AOI2BB1X1TF U907 ( .A0N(N294), .A1N(X_IN[6]), .B0(Y_IN[4]), .Y(N292) );
  AOI2BB1X1TF U908 ( .A0N(N298), .A1N(X_IN[8]), .B0(Y_IN[6]), .Y(N296) );
  NAND2X1TF U909 ( .A(N163), .B(N186), .Y(N617) );
  NAND4BX1TF U910 ( .AN(N381), .B(N316), .C(N804), .D(N364), .Y(N725) );
  NAND2X1TF U911 ( .A(N839), .B(N162), .Y(N847) );
  NAND2X1TF U912 ( .A(N858), .B(N181), .Y(N867) );
  NOR2BX1TF U913 ( .AN(N892), .B(OPER_B[7]), .Y(N895) );
  NAND2X1TF U914 ( .A(N895), .B(N165), .Y(N908) );
  NAND2X1TF U915 ( .A(N923), .B(N166), .Y(N936) );
  NAND2X1TF U916 ( .A(N343), .B(N180), .Y(N348) );
  NAND2X1TF U917 ( .A(N907), .B(N74), .Y(N958) );
  NAND2X1TF U918 ( .A(N566), .B(N958), .Y(N939) );
  NAND2X1TF U919 ( .A(N967), .B(N379), .Y(N574) );
  NAND3X1TF U920 ( .A(N92), .B(N91), .C(N90), .Y(N592) );
  NOR2BX1TF U921 ( .AN(N574), .B(N606), .Y(N571) );
  NAND2X1TF U922 ( .A(PRE_WORK), .B(N354), .Y(N953) );
  NAND2X1TF U923 ( .A(N606), .B(N824), .Y(N347) );
  NAND2X1TF U924 ( .A(N223), .B(N959), .Y(N366) );
  NAND3X1TF U925 ( .A(SIGN_Y), .B(N74), .C(N906), .Y(N825) );
  NAND2X1TF U926 ( .A(N862), .B(N855), .Y(N868) );
  NAND2X1TF U927 ( .A(N881), .B(N882), .Y(N893) );
  NAND2X1TF U928 ( .A(N897), .B(N898), .Y(N909) );
  NAND2X1TF U929 ( .A(N915), .B(N917), .Y(N933) );
  NAND3X1TF U930 ( .A(N606), .B(N603), .C(N168), .Y(N601) );
  NAND2X1TF U931 ( .A(N414), .B(N413), .Y(N422) );
  NAND2X1TF U932 ( .A(N433), .B(N432), .Y(N443) );
  NAND2X1TF U933 ( .A(N453), .B(N452), .Y(N462) );
  NAND2X1TF U934 ( .A(N499), .B(N498), .Y(N1014) );
  AOI222XLTF U935 ( .A0(XTEMP[11]), .A1(N139), .B0(XTEMP[11]), .B1(N497), .C0(
        N139), .C1(N497), .Y(N355) );
  XOR2X1TF U936 ( .A(X_IN[12]), .B(N355), .Y(N360) );
  NAND3X1TF U937 ( .A(N567), .B(POST_WORK), .C(N603), .Y(N376) );
  NAND3BX1TF U938 ( .AN(N366), .B(N949), .C(N967), .Y(N599) );
  NAND3X1TF U939 ( .A(N610), .B(N367), .C(N599), .Y(N943) );
  NAND2X1TF U940 ( .A(N119), .B(N393), .Y(N380) );
  NAND3X1TF U941 ( .A(N383), .B(N122), .C(DP_OP_333_124_4748_N57), .Y(N639) );
  NOR2BX1TF U942 ( .AN(N635), .B(N944), .Y(N543) );
  NAND2X1TF U943 ( .A(N800), .B(SUM_AB[8]), .Y(N424) );
  NAND4X1TF U944 ( .A(N427), .B(N426), .C(N425), .D(N424), .Y(N428) );
  NAND4X1TF U945 ( .A(N438), .B(N437), .C(N436), .D(N435), .Y(N439) );
  NAND4X1TF U946 ( .A(N448), .B(N447), .C(N446), .D(N445), .Y(N449) );
  OAI2BB1X1TF U947 ( .A0N(DIVISION_HEAD[10]), .A1N(N471), .B0(N451), .Y(N713)
         );
  AOI2BB2X1TF U948 ( .B0(X_IN[9]), .B1(N478), .A0N(N478), .A1N(X_IN[9]), .Y(
        N483) );
  NAND3X1TF U949 ( .A(N126), .B(N529), .C(N483), .Y(N479) );
  AOI2BB1X1TF U950 ( .A0N(N509), .A1N(N483), .B0(N513), .Y(N484) );
  AOI2BB2X1TF U951 ( .B0(N487), .B1(N502), .A0N(N502), .A1N(N487), .Y(N494) );
  AOI2BB1X1TF U952 ( .A0N(N509), .A1N(N494), .B0(N513), .Y(N495) );
  AOI2BB2X1TF U953 ( .B0(N139), .B1(N497), .A0N(N497), .A1N(N139), .Y(N510) );
  OAI2BB2XLTF U954 ( .B0(N502), .B1(N609), .A0N(XTEMP[12]), .A1N(N95), .Y(N503) );
  AOI2BB1X1TF U955 ( .A0N(N509), .A1N(N510), .B0(N513), .Y(N511) );
  AOI2BB1X1TF U956 ( .A0N(DIVISION_REMA[2]), .A1N(N518), .B0(DIVISION_HEAD[6]), 
        .Y(N516) );
  OA21XLTF U957 ( .A0(N157), .A1(DIVISION_REMA[4]), .B0(N520), .Y(N522) );
  OA21XLTF U958 ( .A0(N160), .A1(DIVISION_REMA[6]), .B0(N524), .Y(N526) );
  OA21XLTF U959 ( .A0(XTEMP[12]), .A1(N536), .B0(N649), .Y(N535) );
  NAND4X1TF U960 ( .A(N546), .B(N545), .C(N639), .D(N544), .Y(N557) );
  NAND3X1TF U961 ( .A(N552), .B(N551), .C(N550), .Y(N553) );
  NAND3X1TF U962 ( .A(N757), .B(N560), .C(N559), .Y(N561) );
  NAND3X1TF U963 ( .A(N567), .B(N603), .C(N823), .Y(N573) );
  NAND4X1TF U964 ( .A(N569), .B(N568), .C(N640), .D(N573), .Y(N570) );
  NAND2X1TF U965 ( .A(N185), .B(N164), .Y(N591) );
  NOR4XLTF U966 ( .A(\RSHT_BITS[3] ), .B(N90), .C(N615), .D(N591), .Y(N572) );
  NAND2X1TF U967 ( .A(N580), .B(N590), .Y(N587) );
  NAND2X1TF U968 ( .A(N92), .B(N91), .Y(N589) );
  AOI2BB2X1TF U969 ( .B0(N597), .B1(N164), .A0N(N591), .A1N(N593), .Y(N585) );
  NAND4X1TF U970 ( .A(N100), .B(N635), .C(N634), .D(N633), .Y(N636) );
  NAND4X1TF U971 ( .A(N641), .B(N640), .C(N639), .D(N644), .Y(N697) );
  NAND3X1TF U972 ( .A(N757), .B(N653), .C(N652), .Y(N654) );
  AO22X1TF U973 ( .A0(DIVISION_REMA[4]), .A1(N736), .B0(N197), .B1(N791), .Y(
        N744) );
  AOI2BB1X1TF U974 ( .A0N(X_IN[1]), .A1N(N765), .B0(N764), .Y(N768) );
  NAND4X1TF U975 ( .A(N795), .B(N794), .C(N793), .D(N792), .Y(N796) );
  OAI221XLTF U976 ( .A0(\INDEX[2] ), .A1(N90), .B0(N124), .B1(\RSHT_BITS[3] ), 
        .C0(N818), .Y(N819) );
  OAI221XLTF U977 ( .A0(N129), .A1(N185), .B0(N163), .B1(N92), .C0(N820), .Y(
        N836) );
  NAND2X1TF U978 ( .A(N904), .B(N876), .Y(N871) );
  NAND2BX1TF U979 ( .AN(N821), .B(N871), .Y(N891) );
  NAND2X1TF U980 ( .A(N835), .B(N967), .Y(N877) );
  NAND3X1TF U981 ( .A(SIGN_Y), .B(N74), .C(N225), .Y(N843) );
  OAI2BB1X1TF U982 ( .A0N(N960), .A1N(N836), .B0(N835), .Y(N920) );
  NAND3X1TF U983 ( .A(N74), .B(N182), .C(N61), .Y(N975) );
  NAND4X1TF U984 ( .A(N225), .B(N182), .C(N61), .D(N965), .Y(N845) );
  NAND2X1TF U985 ( .A(N904), .B(N920), .Y(N938) );
  NAND2X1TF U986 ( .A(N941), .B(N946), .Y(N947) );
  NAND2X1TF U987 ( .A(N979), .B(N978), .Y(N668) );
  NAND2X1TF U988 ( .A(N982), .B(N981), .Y(N667) );
  NAND2X1TF U989 ( .A(SUM_AB[3]), .B(N88), .Y(N983) );
  NAND2X1TF U990 ( .A(N988), .B(N987), .Y(N665) );
  NAND2X1TF U991 ( .A(SUM_AB[5]), .B(N88), .Y(N989) );
  NAND2X1TF U992 ( .A(N994), .B(N993), .Y(N663) );
  NAND2X1TF U993 ( .A(SUM_AB[7]), .B(N88), .Y(N995) );
  NAND2X1TF U994 ( .A(N1000), .B(N999), .Y(N661) );
  NAND2X1TF U995 ( .A(SUM_AB[9]), .B(N88), .Y(N1001) );
  NAND2X1TF U996 ( .A(N1006), .B(N1005), .Y(N659) );
  NAND2X1TF U997 ( .A(SUM_AB[11]), .B(N88), .Y(N1007) );
endmodule


module SERIAL_CPU_8BIT_VG ( CLK, ENABLE, RST_N, START, I_DATAIN, D_DATAIN, 
        CPU_WAIT, IS_I_ADDR, NXT, I_ADDR, D_ADDR, D_WE, D_DATAOUT, IO_STATUS, 
        IO_DATAINA, IO_DATAINB, IO_DATAOUTA, IO_DATAOUTB, IO_OFFSET, I_PC, 
        I_REG_C, \IO_CONTROL[15] , \IO_CONTROL[14] , \IO_CONTROL[13] , 
        \IO_CONTROL[12] , \IO_CONTROL[11] , \IO_CONTROL[10] , \IO_CONTROL[9] , 
        \IO_CONTROL[8] , \IO_CONTROL[7] , \IO_CONTROL[6] , \IO_CONTROL[5]_BAR , 
        \IO_CONTROL[4] , \IO_CONTROL[3] , \IO_CONTROL[2] , \IO_CONTROL[1] , 
        \IO_CONTROL[0]  );
  input [7:0] I_DATAIN;
  input [7:0] D_DATAIN;
  output [1:0] NXT;
  output [9:0] I_ADDR;
  output [9:0] D_ADDR;
  output [7:0] D_DATAOUT;
  input [15:0] IO_STATUS;
  input [15:0] IO_DATAINA;
  input [15:0] IO_DATAINB;
  output [15:0] IO_DATAOUTA;
  output [15:0] IO_DATAOUTB;
  output [15:0] IO_OFFSET;
  output [5:0] I_PC;
  output [5:0] I_REG_C;
  input CLK, ENABLE, RST_N, START, CPU_WAIT;
  output IS_I_ADDR, D_WE, \IO_CONTROL[15] , \IO_CONTROL[14] , \IO_CONTROL[13] ,
         \IO_CONTROL[12] , \IO_CONTROL[11] , \IO_CONTROL[10] , \IO_CONTROL[9] ,
         \IO_CONTROL[8] , \IO_CONTROL[7] , \IO_CONTROL[6] ,
         \IO_CONTROL[5]_BAR , \IO_CONTROL[4] , \IO_CONTROL[3] ,
         \IO_CONTROL[2] , \IO_CONTROL[1] , \IO_CONTROL[0] ;
  wire   N89, N90, N91, N92, N93, N94, N95, N96, N97, N1375, N1376, N1377,
         N1378, N1379, N1380, N1381, N1382, \IO_CONTROL[5] , N1383, N1384,
         N1385, N1386, N1387, N1388, N1389, N1390, N1391, N1392, N1393, N1394,
         \GR[7][15] , \GR[7][14] , \GR[7][13] , \GR[7][12] , \GR[7][11] ,
         \GR[7][10] , \GR[7][9] , \GR[7][8] , \GR[7][7] , \GR[7][6] ,
         \GR[7][5] , \GR[7][4] , \GR[7][3] , \GR[7][2] , \GR[7][1] ,
         \GR[7][0] , \GR[6][15] , \GR[6][14] , \GR[6][13] , \GR[6][12] ,
         \GR[6][11] , \GR[6][10] , \GR[6][9] , \GR[6][8] , \GR[6][7] ,
         \GR[6][6] , \GR[6][5] , \GR[6][4] , \GR[6][3] , \GR[6][2] ,
         \GR[6][1] , \GR[6][0] , \GR[5][15] , \GR[5][14] , \GR[5][13] ,
         \GR[5][12] , \GR[5][11] , \GR[5][10] , \GR[5][9] , \GR[5][8] ,
         \GR[5][7] , \GR[5][6] , \GR[5][5] , \GR[5][4] , \GR[5][3] ,
         \GR[5][2] , \GR[5][1] , \GR[5][0] , \GR[0][15] , \GR[0][14] ,
         \GR[0][13] , \GR[0][12] , \GR[0][11] , \GR[0][10] , \GR[0][9] ,
         \GR[0][8] , \GR[0][7] , \GR[0][6] , \GR[0][5] , \GR[0][4] ,
         \GR[0][3] , \GR[0][2] , \GR[0][1] , \GR[0][0] , INSTR_OVER, N165,
         N166, N167, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N207, N208, N209, N210,
         N211, N212, N213, N214, N215, N216, N217, N218, N219, N220, N221,
         N222, N247, N248, N249, N250, N251, N252, N253, N254, N255, N256,
         N257, N258, N259, N260, N261, N262, CF_BUF, N457, N458, N459, N460,
         N461, N462, N463, N464, N465, N466, N467, N468, N469, N470, N471,
         N472, N473, N491, N492, N493, N494, N495, N496, N497, N498, N499,
         N500, N501, N502, N503, N504, N505, N506, N575, N576, ZF, NF, CF,
         N603, N882, N2540, N2550, N2560, N2570, N2580, N2590, N2600, N2610,
         N2620, N287, N288, N289, N293, N294, N295, N296, N297, N298, N299,
         N300, N301, N302, N303, N304, N305, N306, N307, N308, N318, N328,
         N338, N348, N358, N368, N378, N388, N398, N408, N418, N428, N438,
         N448, N4580, N4680, N4690, N4700, N4710, N4720, N4730, N474, N475,
         N476, N477, N478, N479, N480, N481, N482, N483, N484, N485, N486,
         N487, N488, N489, N490, N4910, N4920, N4930, N4940, N4950, N4960,
         N4970, N4980, N4990, N5000, N5010, N5020, N5030, N5040, N5050, N5060,
         N507, N508, N513, N515, N516, N517, N518, N519, N520, N545, N546,
         N560, N565, N566, N567, N568, N569, N570, N571, N572, N573, N574,
         N5750, N5760, N599, N713, N717, N718, N719, N720, N721, N722, N775,
         N776, N831, N832, N833, N834, N835, N836, N837, N838, N839, N840,
         N841, N842, N843, N844, N845, N846, N847, N848, N849, N850, N851,
         N852, N853, N854, N855, N856, N857, N858, N859, N860, N861, N862,
         N863, N864, N865, N866, N867, N868, N869, N870, N871, N872, N873,
         N874, N875, N876, N877, N878, N879, N880, N881, N8820, N883, N884,
         N885, N886, N887, N888, N889, N890, N891, N892, N893, N894, N895,
         N896, N897, N898, N899, N900, N901, N902, N903, N904, N905, N906,
         N907, N908, N909, N910, N911, N912, N913, N914, N915, N916, N917,
         N918, N919, N920, N921, N922, N923, N924, N925, N926, N927, N928,
         N929, N930, N931, N932, N933, N934, N935, N936, N937, N938, N939,
         N940, N941, N942, N943, N944, N945, N946, N947, N948, N949, N950,
         N951, N952, N953, N954, N955, N956, N957, N958, N959, N960,
         ADD_X_299_3_N22, ADD_X_299_3_N21, ADD_X_299_3_N20, ADD_X_299_3_N19,
         ADD_X_299_3_N18, ADD_X_299_3_N17, ADD_X_299_3_N16, ADD_X_299_3_N15,
         ADD_X_299_3_N14, ADD_X_299_3_N13, ADD_X_299_3_N12, ADD_X_299_3_N11,
         ADD_X_299_3_N10, ADD_X_299_3_N9, ADD_X_299_3_N8, ADD_X_299_3_N7,
         ADD_X_299_3_N6, ADD_X_299_3_N5, ADD_X_299_3_N4, ADD_X_299_3_N3,
         ADD_X_299_3_N2, SUB_X_299_4_N16, SUB_X_299_4_N15, SUB_X_299_4_N14,
         SUB_X_299_4_N13, SUB_X_299_4_N12, SUB_X_299_4_N11, SUB_X_299_4_N10,
         SUB_X_299_4_N9, SUB_X_299_4_N8, SUB_X_299_4_N7, SUB_X_299_4_N6,
         SUB_X_299_4_N5, SUB_X_299_4_N4, SUB_X_299_4_N3, SUB_X_299_4_N2,
         SUB_X_299_4_N1, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12,
         N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26,
         N27, N28, N29, N30, N31, N32, N33, N34, N35, N1700, N188, N189, N191,
         N193, N195, N197, N198, N199, N200, N201, N202, N204, N206, N2080,
         N2100, N2110, N2130, N2140, N2150, N2160, N2170, N2190, N2200, N2210,
         N2220, N223, N224, N225, N226, N227, N228, N229, N230, N231, N232,
         N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243,
         N244, N245, N246, N2470, N2480, N2490, N2500, N2510, N2520, N2530,
         N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, N273,
         N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284,
         N285, N286, N290, N291, N292, N309, N310, N311, N312, N313, N314,
         N315, N316, N317, N319, N320, N321, N323, N325, N326, N327, N330,
         N331, N332, N333, N334, N335, N336, N337, N339, N340, N341, N342,
         N343, N344, N345, N346, N347, N349, N350, N351, N352, N370, N371,
         N372, N373, N374, N375, N376, N377, N379, N380, N381, N382, N383,
         N384, N385, N386, N387, N389, N390, N391, N392, N393, N394, N395,
         N396, N397, N399, N400, N401, N402, N403, N404, N405, N406, N407,
         N409, N410, N411, N412, N413, N414, N415, N416, N417, N419, N420,
         N421, N422, N423, N424, N425, N426, N427, N429, N430, N431, N432,
         N433, N434, N435, N436, N437, N439, N440, N441, N442, N443, N444,
         N445, N446, N447, N449, N450, N451, N452, N453, N454, N455, N456,
         N4570, N4590, N4600, N4610, N4620, N4630, N4640, N4650, N4660, N4670,
         N510, N511, N512, N514, N521, N522, N523, N524, N525, N526, N527,
         N528, N529, N530, N531, N532, N533, N534, N535, N536, N537, N538,
         N539, N540, N541, N542, N543, N544, N547, N548, N549, N550, N551,
         N552, N553, N554, N555, N556, N557, N558, N559, N561, N562, N563,
         N564, N577, N578, N579, N580, N581, N582, N583, N584, N585, N586,
         N587, N588, N589, N590, N591, N592, N593, N594, N595, N596, N597,
         N598, N600, N601, N602, N6030, N604, N605, N606, N607, N608, N609,
         N610, N611, N612, N613, N614, N615, N616, N617, N618, N619, N620,
         N621, N622, N623, N624, N625, N626, N627, N628, N629, N630, N631,
         N632, N633, N634, N635, N636, N637, N638, N639, N640, N641, N642,
         N643, N644, N645, N646, N647, N648, N649, N650, N651, N652, N653,
         N654, N655, N656, N657, N658, N659, N660, N661, N662, N663, N664,
         N665, N666, N667, N668, N669, N670, N671, N672, N673, N674, N675,
         N676, N677, N678, N679, N680, N681, N682, N683, N684, N685, N686,
         N687, N688, N689, N690, N691, N692, N693, N694, N695, N696, N697,
         N698, N699, N700, N701, N702, N703, N704, N705, N706, N707, N708,
         N709, N710, N711, N712, N714, N715, N716, N723, N724, N725, N726,
         N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737,
         N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748,
         N749, N750, N751, N752, N753, N754, N755, N756, N757, N758, N759,
         N760, N761, N762, N763, N764, N765, N766, N767, N768, N769, N770,
         N771, N772, N773, N774, N777, N778, N779, N780, N781, N782, N783,
         N784, N785, N786, N787, N788, N789, N790, N791, N792, N793, N794,
         N795, N796, N797, N798, N799, N800, N801, N802, N803, N804, N805,
         N806, N807, N808, N809, N810, N811, N812, N813, N814, N815, N816,
         N817, N818, N819, N820, N821, N822, N823, N824, N825, N826, N827,
         N828, N829, N830, N961, N962, N963, N964, N965, N966, N967, N968,
         N969, N970, N971, N972, N973, N974, N975, N976, N977, N978, N979,
         N980, N981, N982, N983, N984, N985, N986, N987, N988, N989, N990,
         N991, N992, N993, N994, N995, N996, N997, N998, N999, N1000, N1001,
         N1002, N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011,
         N1012, N1013, N1014, N1015, N1016, N1017, N1018, N1019, N1020, N1021,
         N1022, N1023, N1024, N1025, N1026, N1027, N1028, N1029, N1030, N1031,
         N1032, N1033, N1034, N1035, N1036, N1037, N1038, N1039, N1040, N1041,
         N1042, N1043, N1044, N1045, N1046, N1047, N1048, N1049, N1050, N1051,
         N1052, N1053, N1054, N1055, N1056, N1057, N1058, N1059, N1060, N1061,
         N1062, N1063, N1064, N1065, N1066, N1067, N1068, N1069, N1070, N1071,
         N1072, N1073, N1074, N1075, N1076, N1077, N1078, N1079, N1080, N1081,
         N1082, N1083, N1084, N1085, N1086, N1087, N1088, N1089, N1090, N1091,
         N1092, N1093, N1094, N1095, N1096, N1097, N1098, N1099, N1100, N1101,
         N1102, N1103, N1104, N1105, N1106, N1107, N1108, N1109, N1110, N1111,
         N1112, N1113, N1114, N1115, N1116, N1117, N1118, N1119, N1120, N1121,
         N1122, N1123, N1124, N1125, N1126, N1127, N1128, N1129, N1130, N1131,
         N1132, N1133, N1134, N1135, N1136, N1137, N1138, N1139, N1140, N1141,
         N1142, N1143, N1144, N1145, N1146, N1147, N1148, N1149, N1150, N1151,
         N1152, N1153, N1154, N1155, N1156, N1157, N1158, N1159, N1160, N1161,
         N1162, N1163, N1164, N1165, N1166, N1167, N1168, N1169, N1170, N1171,
         N1172, N1173, N1174, N1175, N1176, N1177, N1178, N1179, N1180, N1181,
         N1182, N1183, N1184, N1185, N1186, N1187, N1188, N1189, N1190, N1191,
         N1192, N1193, N1194, N1195, N1196, N1197, N1198, N1199, N1200, N1201,
         N1202, N1203, N1204, N1205, N1206, N1207, N1208, N1209, N1210, N1211,
         N1212, N1213, N1214, N1215, N1216, N1217, N1218, N1219, N1220, N1221,
         N1222, N1223, N1224, N1225, N1226, N1227, N1228, N1229, N1230, N1231,
         N1232, N1233, N1234, N1235, N1236, N1237, N1238, N1239, N1240, N1241,
         N1242, N1243, N1244, N1245, N1246, N1247, N1248, N1249, N1250, N1251,
         N1252, N1253, N1254, N1255, N1256, N1257, N1258, N1259, N1260, N1261,
         N1262, N1263, N1264, N1265, N1266, N1267, N1268, N1269, N1270, N1271,
         N1272, N1273, N1274, N1275, N1276, N1277, N1278, N1279, N1280, N1281,
         N1282, N1283, N1284, N1285, N1286, N1287, N1288, N1289, N1290, N1291,
         N1292, N1293, N1294, N1295, N1296, N1297, N1298, N1299, N1300, N1301,
         N1302, N1303, N1304, N1305, N1306, N1307, N1308, N1309, N1310, N1311,
         N1312, N1313, N1314, N1315, N1316, N1317, N1318, N1319, N1320, N1321,
         N1322, N1323, N1324, N1325, N1326, N1327, N1328, N1329, N1330, N1331,
         N1332, N1333, N1334, N1335, N1336, N1337, N1338, N1339, N1340, N1341,
         N1342, N1343, N1344, N1345, N1346, N1347, N1348, N1349, N1350, N1351,
         N1352, N1353, N1354, N1355, N1356, N1357, N1358, N1359, N1360, N1361,
         N1362, N1363, N1364, N1365, N1366, N1367, N1368, N1369, N1370, N1371,
         N1372, N1373, N1374;
  wire   [3:1] CODE_TYPE;
  wire   [3:1] STATE;
  wire   [3:0] NEXT_STATE;
  wire   [15:0] REG_A;
  wire   [15:0] REG_B;
  wire   [15:0] SMDR;

  DFFRX4TF \reg_B_reg[0]  ( .D(N485), .CK(CLK), .RN(RST_N), .Q(REG_B[0]), .QN(
        N371) );
  CLKINVX6TF U404 ( .A(RST_N), .Y(N599) );
  AFCSIHCONX2TF \add_x_299_3/U17  ( .A(REG_B[2]), .B(REG_A[2]), .CS(
        ADD_X_299_3_N21), .S(N459), .CO0N(ADD_X_299_3_N20), .CO1N(
        ADD_X_299_3_N19) );
  AFCSHCINX2TF \add_x_299_3/U16  ( .CI1N(ADD_X_299_3_N19), .B(REG_B[3]), .A(
        REG_A[3]), .CI0N(ADD_X_299_3_N20), .CS(ADD_X_299_3_N21), .CO1(
        ADD_X_299_3_N17), .CO0(ADD_X_299_3_N18), .S(N460) );
  AFCSIHCONX2TF \add_x_299_3/U14  ( .A(REG_A[4]), .B(REG_B[4]), .CS(
        ADD_X_299_3_N16), .S(N461), .CO0N(ADD_X_299_3_N15), .CO1N(
        ADD_X_299_3_N14) );
  AFCSHCINX2TF \add_x_299_3/U13  ( .CI1N(ADD_X_299_3_N14), .B(REG_A[5]), .A(
        REG_B[5]), .CI0N(ADD_X_299_3_N15), .CS(ADD_X_299_3_N16), .CO1(
        ADD_X_299_3_N12), .CO0(ADD_X_299_3_N13), .S(N462) );
  CMPR32X2TF \add_x_299_3/U11  ( .A(REG_A[6]), .B(REG_B[6]), .C(
        ADD_X_299_3_N11), .CO(ADD_X_299_3_N10), .S(N463) );
  CMPR32X2TF \add_x_299_3/U10  ( .A(REG_A[7]), .B(REG_B[7]), .C(
        ADD_X_299_3_N10), .CO(ADD_X_299_3_N9), .S(N464) );
  CMPR32X2TF \add_x_299_3/U9  ( .A(REG_A[8]), .B(REG_B[8]), .C(ADD_X_299_3_N9), 
        .CO(ADD_X_299_3_N8), .S(N465) );
  CMPR32X2TF \add_x_299_3/U8  ( .A(REG_A[9]), .B(REG_B[9]), .C(ADD_X_299_3_N8), 
        .CO(ADD_X_299_3_N7), .S(N466) );
  CMPR32X2TF \add_x_299_3/U7  ( .A(REG_A[10]), .B(REG_B[10]), .C(
        ADD_X_299_3_N7), .CO(ADD_X_299_3_N6), .S(N467) );
  CMPR32X2TF \add_x_299_3/U6  ( .A(REG_A[11]), .B(REG_B[11]), .C(
        ADD_X_299_3_N6), .CO(ADD_X_299_3_N5), .S(N468) );
  CMPR32X2TF \add_x_299_3/U5  ( .A(REG_A[12]), .B(REG_B[12]), .C(
        ADD_X_299_3_N5), .CO(ADD_X_299_3_N4), .S(N469) );
  CMPR32X2TF \add_x_299_3/U4  ( .A(REG_A[13]), .B(REG_B[13]), .C(
        ADD_X_299_3_N4), .CO(ADD_X_299_3_N3), .S(N470) );
  CMPR32X2TF \add_x_299_3/U3  ( .A(REG_A[14]), .B(REG_B[14]), .C(
        ADD_X_299_3_N3), .CO(ADD_X_299_3_N2), .S(N471) );
  DFFSX2TF \pc_reg[7]  ( .D(N713), .CK(CLK), .SN(RST_N), .Q(N423), .QN(
        I_ADDR[8]) );
  DFFSX2TF \pc_reg[3]  ( .D(N720), .CK(CLK), .SN(RST_N), .Q(N422), .QN(
        I_ADDR[4]) );
  DFFSX2TF \pc_reg[1]  ( .D(N722), .CK(CLK), .SN(RST_N), .Q(N421), .QN(
        I_ADDR[2]) );
  DFFSX2TF \pc_reg[5]  ( .D(N718), .CK(CLK), .SN(RST_N), .Q(N420), .QN(
        I_ADDR[6]) );
  DFFSX2TF \pc_reg[0]  ( .D(N776), .CK(CLK), .SN(RST_N), .Q(N419), .QN(
        I_ADDR[1]) );
  DFFSX2TF \pc_reg[8]  ( .D(N775), .CK(CLK), .SN(RST_N), .Q(N417), .QN(
        I_ADDR[9]) );
  DFFRX2TF nf_reg ( .D(N288), .CK(CLK), .RN(RST_N), .Q(NF), .QN(N416) );
  DFFSX2TF \pc_reg[6]  ( .D(N717), .CK(CLK), .SN(RST_N), .Q(N415), .QN(
        I_ADDR[7]) );
  DFFSX2TF \pc_reg[4]  ( .D(N719), .CK(CLK), .SN(RST_N), .Q(N414), .QN(
        I_ADDR[5]) );
  DFFSX2TF \pc_reg[2]  ( .D(N721), .CK(CLK), .SN(RST_N), .Q(N413), .QN(
        I_ADDR[3]) );
  DFFRX2TF \reg_B_reg[10]  ( .D(N4950), .CK(CLK), .RN(RST_N), .Q(REG_B[10]), 
        .QN(N570) );
  DFFRX2TF \reg_A_reg[10]  ( .D(N479), .CK(CLK), .RN(RST_N), .Q(REG_A[10]), 
        .QN(N411) );
  DFFRX2TF \reg_A_reg[11]  ( .D(N480), .CK(CLK), .RN(RST_N), .Q(REG_A[11]), 
        .QN(N410) );
  DFFRX2TF \state_reg[2]  ( .D(NEXT_STATE[2]), .CK(CLK), .RN(RST_N), .Q(N409), 
        .QN(N545) );
  DFFRX2TF \reg_B_reg[3]  ( .D(N488), .CK(CLK), .RN(RST_N), .Q(REG_B[3]), .QN(
        N407) );
  DFFRX2TF \reg_B_reg[1]  ( .D(N486), .CK(CLK), .RN(RST_N), .Q(REG_B[1]), .QN(
        N406) );
  DFFRX2TF \reg_B_reg[2]  ( .D(N487), .CK(CLK), .RN(RST_N), .Q(REG_B[2]), .QN(
        N405) );
  DFFRX2TF \id_ir_reg[1]  ( .D(N507), .CK(CLK), .RN(RST_N), .Q(N96), .QN(N404)
         );
  DFFRX2TF \id_ir_reg[5]  ( .D(N5030), .CK(CLK), .RN(RST_N), .Q(N93), .QN(N403) );
  DFFRX2TF \reg_A_reg[12]  ( .D(N481), .CK(CLK), .RN(RST_N), .Q(REG_A[12]), 
        .QN(N402) );
  DFFRX2TF \reg_A_reg[13]  ( .D(N482), .CK(CLK), .RN(RST_N), .Q(REG_A[13]), 
        .QN(N401) );
  DFFRX2TF \reg_A_reg[8]  ( .D(N477), .CK(CLK), .RN(RST_N), .Q(REG_A[8]), .QN(
        N400) );
  DFFRX2TF \reg_A_reg[7]  ( .D(N476), .CK(CLK), .RN(RST_N), .Q(REG_A[7]), .QN(
        N399) );
  DFFRX2TF \reg_A_reg[9]  ( .D(N478), .CK(CLK), .RN(RST_N), .Q(REG_A[9]), .QN(
        N397) );
  DFFRX2TF \reg_A_reg[6]  ( .D(N475), .CK(CLK), .RN(RST_N), .Q(REG_A[6]), .QN(
        N396) );
  DFFRX2TF \state_reg[1]  ( .D(NEXT_STATE[1]), .CK(CLK), .RN(RST_N), .Q(
        STATE[1]), .QN(N395) );
  DFFRX2TF \reg_A_reg[2]  ( .D(N4710), .CK(CLK), .RN(RST_N), .Q(REG_A[2]), 
        .QN(N394) );
  DFFRX2TF \reg_A_reg[4]  ( .D(N4730), .CK(CLK), .RN(RST_N), .Q(REG_A[4]), 
        .QN(N393) );
  DFFRX2TF \reg_A_reg[15]  ( .D(N484), .CK(CLK), .RN(RST_N), .Q(REG_A[15]), 
        .QN(N391) );
  DFFRX2TF \id_ir_reg[13]  ( .D(N515), .CK(CLK), .RN(RST_N), .Q(CODE_TYPE[2]), 
        .QN(N390) );
  DFFRX2TF \reg_A_reg[3]  ( .D(N4720), .CK(CLK), .RN(RST_N), .Q(REG_A[3]), 
        .QN(N389) );
  DFFRX2TF \reg_A_reg[5]  ( .D(N474), .CK(CLK), .RN(RST_N), .Q(REG_A[5]), .QN(
        N387) );
  DFFRX2TF \reg_A_reg[1]  ( .D(N4700), .CK(CLK), .RN(RST_N), .Q(REG_A[1]), 
        .QN(N386) );
  DFFRX2TF \id_ir_reg[15]  ( .D(N513), .CK(CLK), .RN(RST_N), .Q(N22), .QN(N384) );
  DFFRX2TF \id_ir_reg[0]  ( .D(N508), .CK(CLK), .RN(RST_N), .Q(N95), .QN(N383)
         );
  DFFRX2TF \id_ir_reg[4]  ( .D(N5040), .CK(CLK), .RN(RST_N), .Q(N92), .QN(N382) );
  DFFRX2TF \id_ir_reg[8]  ( .D(N520), .CK(CLK), .RN(RST_N), .Q(N89), .QN(N381)
         );
  DFFRX2TF \id_ir_reg[9]  ( .D(N519), .CK(CLK), .RN(RST_N), .Q(N90), .QN(N380)
         );
  DFFRX2TF \reg_A_reg[14]  ( .D(N483), .CK(CLK), .RN(RST_N), .Q(REG_A[14]), 
        .QN(N379) );
  DFFRX2TF \id_ir_reg[6]  ( .D(N5020), .CK(CLK), .RN(RST_N), .Q(N94), .QN(N376) );
  DFFRX2TF \id_ir_reg[2]  ( .D(N5060), .CK(CLK), .RN(RST_N), .Q(N97), .QN(N375) );
  DFFRX2TF \id_ir_reg[10]  ( .D(N518), .CK(CLK), .RN(RST_N), .Q(N91), .QN(N374) );
  DFFRX2TF \state_reg[0]  ( .D(NEXT_STATE[0]), .CK(CLK), .RN(RST_N), .Q(N370), 
        .QN(N546) );
  TLATXLTF cf_buf_reg ( .G(N575), .D(N576), .Q(CF_BUF) );
  TLATXLTF \nxt_reg[1]  ( .G(N165), .D(N167), .Q(NXT[1]) );
  TLATXLTF \nxt_reg[0]  ( .G(N165), .D(N166), .Q(NXT[0]) );
  DFFRX2TF \id_ir_reg[7]  ( .D(N5010), .CK(CLK), .RN(RST_N), .QN(N2550) );
  DFFRX2TF \id_ir_reg[3]  ( .D(N5050), .CK(CLK), .RN(RST_N), .QN(N2540) );
  DFFRX2TF \reg_B_reg[15]  ( .D(N5000), .CK(CLK), .RN(RST_N), .Q(REG_B[15]), 
        .QN(N565) );
  DFFRX2TF \reg_B_reg[14]  ( .D(N4990), .CK(CLK), .RN(RST_N), .Q(REG_B[14]), 
        .QN(N566) );
  DFFRX2TF \reg_B_reg[13]  ( .D(N4980), .CK(CLK), .RN(RST_N), .Q(REG_B[13]), 
        .QN(N567) );
  DFFRX2TF \reg_B_reg[12]  ( .D(N4970), .CK(CLK), .RN(RST_N), .Q(REG_B[12]), 
        .QN(N568) );
  DFFRX2TF \reg_B_reg[11]  ( .D(N4960), .CK(CLK), .RN(RST_N), .Q(REG_B[11]), 
        .QN(N569) );
  DFFNSRX2TF is_i_addr_reg ( .D(N959), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        IS_I_ADDR) );
  DFFNSRX2TF \reg_C_reg[7]  ( .D(N4680), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[8]) );
  DFFNSRX2TF \reg_C_reg[6]  ( .D(N4580), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[7]) );
  DFFNSRX2TF \reg_C_reg[8]  ( .D(N338), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[9]) );
  DFFRX2TF \reg_B_reg[9]  ( .D(N4940), .CK(CLK), .RN(RST_N), .Q(REG_B[9]), 
        .QN(N571) );
  DFFRX2TF \reg_B_reg[8]  ( .D(N4930), .CK(CLK), .RN(RST_N), .Q(REG_B[8]), 
        .QN(N572) );
  DFFRX2TF \reg_B_reg[7]  ( .D(N4920), .CK(CLK), .RN(RST_N), .Q(REG_B[7]), 
        .QN(N573) );
  DFFRX2TF \reg_B_reg[6]  ( .D(N4910), .CK(CLK), .RN(RST_N), .Q(REG_B[6]), 
        .QN(N574) );
  DFFRX2TF \reg_B_reg[5]  ( .D(N490), .CK(CLK), .RN(RST_N), .Q(REG_B[5]), .QN(
        N5750) );
  DFFRX2TF \reg_B_reg[4]  ( .D(N489), .CK(CLK), .RN(RST_N), .Q(REG_B[4]), .QN(
        N5760) );
  DFFNSRX2TF \reg_C_reg[5]  ( .D(N388), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[6]) );
  DFFNSRX2TF \reg_C_reg[1]  ( .D(N328), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[2]) );
  DFFNSRX2TF \reg_C_reg[3]  ( .D(N428), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[4]) );
  DFFNSRX2TF \reg_C_reg[4]  ( .D(N378), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[5]) );
  DFFNSRX2TF \reg_C_reg[2]  ( .D(N418), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[3]) );
  DFFNSRX2TF \reg_C_reg[0]  ( .D(N318), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[1]) );
  DFFRX2TF \id_ir_reg[12]  ( .D(N516), .CK(CLK), .RN(RST_N), .Q(CODE_TYPE[1]), 
        .QN(N377) );
  ADDHXLTF \add_x_299_3/U19  ( .A(REG_B[0]), .B(REG_A[0]), .CO(ADD_X_299_3_N22), .S(N457) );
  CMPR32X2TF \add_x_299_3/U2  ( .A(REG_A[15]), .B(REG_B[15]), .C(
        ADD_X_299_3_N2), .CO(N473), .S(N472) );
  CMPR32X2TF \add_x_299_3/U18  ( .A(REG_A[1]), .B(REG_B[1]), .C(
        ADD_X_299_3_N22), .CO(ADD_X_299_3_N21), .S(N458) );
  CLKMX2X2TF \add_x_299_3/U12  ( .A(ADD_X_299_3_N13), .B(ADD_X_299_3_N12), 
        .S0(ADD_X_299_3_N16), .Y(ADD_X_299_3_N11) );
  CLKMX2X4TF \add_x_299_3/U15  ( .A(ADD_X_299_3_N18), .B(ADD_X_299_3_N17), 
        .S0(ADD_X_299_3_N21), .Y(ADD_X_299_3_N16) );
  DFFRX4TF \reg_A_reg[0]  ( .D(N4690), .CK(CLK), .RN(RST_N), .Q(REG_A[0]), 
        .QN(N392) );
  CMPR32X2TF \sub_x_299_4/U6  ( .A(N569), .B(REG_A[11]), .C(SUB_X_299_4_N6), 
        .CO(SUB_X_299_4_N5), .S(N502) );
  CMPR32X2TF \sub_x_299_4/U10  ( .A(N573), .B(REG_A[7]), .C(SUB_X_299_4_N10), 
        .CO(SUB_X_299_4_N9), .S(N498) );
  CMPR32X2TF \sub_x_299_4/U11  ( .A(N574), .B(REG_A[6]), .C(SUB_X_299_4_N11), 
        .CO(SUB_X_299_4_N10), .S(N497) );
  CMPR32X2TF \sub_x_299_4/U12  ( .A(N5750), .B(REG_A[5]), .C(SUB_X_299_4_N12), 
        .CO(SUB_X_299_4_N11), .S(N496) );
  CMPR32X2TF \sub_x_299_4/U9  ( .A(N572), .B(REG_A[8]), .C(SUB_X_299_4_N9), 
        .CO(SUB_X_299_4_N8), .S(N499) );
  CMPR32X2TF \sub_x_299_4/U15  ( .A(N405), .B(REG_A[2]), .C(SUB_X_299_4_N15), 
        .CO(SUB_X_299_4_N14), .S(N493) );
  CMPR32X2TF \sub_x_299_4/U7  ( .A(N570), .B(REG_A[10]), .C(SUB_X_299_4_N7), 
        .CO(SUB_X_299_4_N6), .S(N501) );
  CMPR32X2TF \sub_x_299_4/U5  ( .A(N568), .B(REG_A[12]), .C(SUB_X_299_4_N5), 
        .CO(SUB_X_299_4_N4), .S(N503) );
  INVX2TF \sub_x_299_4/*cell*4322  ( .A(REG_B[3]), .Y(N352) );
  CMPR32X2TF \sub_x_299_4/U3  ( .A(N566), .B(REG_A[14]), .C(SUB_X_299_4_N3), 
        .CO(SUB_X_299_4_N2), .S(N505) );
  CMPR32X2TF \sub_x_299_4/U16  ( .A(N406), .B(REG_A[1]), .C(SUB_X_299_4_N16), 
        .CO(SUB_X_299_4_N15), .S(N492) );
  CMPR32X2TF \sub_x_299_4/U4  ( .A(N567), .B(REG_A[13]), .C(SUB_X_299_4_N4), 
        .CO(SUB_X_299_4_N3), .S(N504) );
  DFFNSRX2TF lowest_bit_reg ( .D(N960), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        I_ADDR[0]), .QN(N412) );
  DFFNSRXLTF \reg_C_reg[10]  ( .D(N408), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N2580) );
  DFFNSRXLTF \reg_C_reg[9]  ( .D(N348), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N2620) );
  DFFNSRXLTF \reg_C_reg[13]  ( .D(N368), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N2600) );
  DFFNSRXLTF \reg_C_reg[12]  ( .D(N358), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N2610) );
  DFFNSRXLTF \reg_C_reg[11]  ( .D(N398), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N2590) );
  DFFNSRXLTF \reg_C_reg[14]  ( .D(N438), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N2570) );
  DFFNSRXLTF \reg_C_reg[15]  ( .D(N448), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N2560) );
  DFFNSRXLTF dw_reg ( .D(N603), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(D_WE) );
  DFFSX2TF \id_ir_reg[14]  ( .D(N1700), .CK(CLK), .SN(RST_N), .Q(N614), .QN(
        CODE_TYPE[3]) );
  DFFRX1TF \state_reg[3]  ( .D(NEXT_STATE[3]), .CK(CLK), .RN(RST_N), .Q(
        STATE[3]), .QN(N752) );
  DFFRX1TF \smdr_reg[15]  ( .D(N308), .CK(CLK), .RN(RST_N), .Q(SMDR[15]) );
  DFFRX1TF \smdr_reg[14]  ( .D(N307), .CK(CLK), .RN(RST_N), .Q(SMDR[14]) );
  DFFRX1TF \smdr_reg[13]  ( .D(N306), .CK(CLK), .RN(RST_N), .Q(SMDR[13]) );
  DFFRX1TF \smdr_reg[6]  ( .D(N299), .CK(CLK), .RN(RST_N), .Q(SMDR[6]) );
  DFFRX1TF \smdr_reg[4]  ( .D(N297), .CK(CLK), .RN(RST_N), .Q(SMDR[4]) );
  DFFRX1TF \smdr_reg[3]  ( .D(N296), .CK(CLK), .RN(RST_N), .Q(SMDR[3]) );
  DFFRX1TF \smdr_reg[2]  ( .D(N295), .CK(CLK), .RN(RST_N), .Q(SMDR[2]) );
  DFFRX1TF \smdr_reg[0]  ( .D(N293), .CK(CLK), .RN(RST_N), .Q(SMDR[0]) );
  DFFRX1TF \smdr_reg[12]  ( .D(N305), .CK(CLK), .RN(RST_N), .Q(SMDR[12]) );
  DFFRX1TF \smdr_reg[11]  ( .D(N304), .CK(CLK), .RN(RST_N), .Q(SMDR[11]) );
  DFFRX1TF \smdr_reg[10]  ( .D(N303), .CK(CLK), .RN(RST_N), .Q(SMDR[10]) );
  DFFRX1TF \smdr_reg[9]  ( .D(N302), .CK(CLK), .RN(RST_N), .Q(SMDR[9]) );
  DFFRX1TF \smdr_reg[8]  ( .D(N301), .CK(CLK), .RN(RST_N), .Q(SMDR[8]) );
  DFFRX1TF \smdr_reg[7]  ( .D(N300), .CK(CLK), .RN(RST_N), .Q(SMDR[7]) );
  DFFRX1TF \smdr_reg[5]  ( .D(N298), .CK(CLK), .RN(RST_N), .Q(SMDR[5]) );
  DFFRX1TF \smdr_reg[1]  ( .D(N294), .CK(CLK), .RN(RST_N), .Q(SMDR[1]) );
  DFFRX1TF cf_reg ( .D(N289), .CK(CLK), .RN(RST_N), .Q(CF) );
  DFFRX1TF instr_over_reg ( .D(N882), .CK(CLK), .RN(RST_N), .Q(INSTR_OVER) );
  DFFRX1TF zf_reg ( .D(N287), .CK(CLK), .RN(RST_N), .Q(ZF) );
  DFFRX1TF \gr_reg[7][12]  ( .D(N834), .CK(CLK), .RN(RST_N), .Q(\GR[7][12] )
         );
  DFFRX1TF \gr_reg[7][11]  ( .D(N835), .CK(CLK), .RN(RST_N), .Q(\GR[7][11] )
         );
  DFFRX1TF \gr_reg[7][10]  ( .D(N836), .CK(CLK), .RN(RST_N), .Q(\GR[7][10] )
         );
  DFFRX1TF \gr_reg[7][9]  ( .D(N837), .CK(CLK), .RN(RST_N), .Q(\GR[7][9] ) );
  DFFRX1TF \gr_reg[6][12]  ( .D(N842), .CK(CLK), .RN(RST_N), .Q(\GR[6][12] )
         );
  DFFRX1TF \gr_reg[6][11]  ( .D(N843), .CK(CLK), .RN(RST_N), .Q(\GR[6][11] )
         );
  DFFRX1TF \gr_reg[6][10]  ( .D(N844), .CK(CLK), .RN(RST_N), .Q(\GR[6][10] )
         );
  DFFRX1TF \gr_reg[6][9]  ( .D(N845), .CK(CLK), .RN(RST_N), .Q(\GR[6][9] ) );
  DFFRX1TF \gr_reg[5][12]  ( .D(N850), .CK(CLK), .RN(RST_N), .Q(\GR[5][12] )
         );
  DFFRX1TF \gr_reg[5][11]  ( .D(N851), .CK(CLK), .RN(RST_N), .Q(\GR[5][11] )
         );
  DFFRX1TF \gr_reg[5][10]  ( .D(N852), .CK(CLK), .RN(RST_N), .Q(\GR[5][10] )
         );
  DFFRX1TF \gr_reg[5][9]  ( .D(N853), .CK(CLK), .RN(RST_N), .Q(\GR[5][9] ) );
  DFFRX1TF \gr_reg[4][12]  ( .D(N858), .CK(CLK), .RN(RST_N), .Q(N1392) );
  DFFRX1TF \gr_reg[4][11]  ( .D(N859), .CK(CLK), .RN(RST_N), .Q(N1393) );
  DFFRX1TF \gr_reg[4][10]  ( .D(N860), .CK(CLK), .RN(RST_N), .Q(N1394) );
  DFFRX1TF \gr_reg[4][9]  ( .D(N861), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[9])
         );
  DFFRX1TF \gr_reg[3][11]  ( .D(N867), .CK(CLK), .RN(RST_N), .Q(N35), .QN(
        N2080) );
  DFFRX1TF \gr_reg[2][12]  ( .D(N874), .CK(CLK), .RN(RST_N), .Q(N34), .QN(N206) );
  DFFRX1TF \gr_reg[2][11]  ( .D(N875), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTA[11]) );
  DFFRX1TF \gr_reg[2][10]  ( .D(N876), .CK(CLK), .RN(RST_N), .Q(N33), .QN(N191) );
  DFFRX1TF \gr_reg[2][9]  ( .D(N877), .CK(CLK), .RN(RST_N), .Q(N32), .QN(N327)
         );
  DFFRX1TF \gr_reg[1][12]  ( .D(N8820), .CK(CLK), .RN(RST_N), .Q(N1378) );
  DFFRX1TF \gr_reg[1][11]  ( .D(N883), .CK(CLK), .RN(RST_N), .Q(N1379) );
  DFFRX1TF \gr_reg[1][10]  ( .D(N884), .CK(CLK), .RN(RST_N), .Q(N1380) );
  DFFRX1TF \gr_reg[1][9]  ( .D(N885), .CK(CLK), .RN(RST_N), .Q(N1381) );
  DFFRX1TF \gr_reg[0][12]  ( .D(N890), .CK(CLK), .RN(RST_N), .Q(\GR[0][12] )
         );
  DFFRX1TF \gr_reg[0][11]  ( .D(N891), .CK(CLK), .RN(RST_N), .Q(\GR[0][11] )
         );
  DFFRX1TF \gr_reg[0][10]  ( .D(N892), .CK(CLK), .RN(RST_N), .Q(\GR[0][10] )
         );
  DFFRX1TF \gr_reg[0][9]  ( .D(N893), .CK(CLK), .RN(RST_N), .Q(\GR[0][9] ) );
  DFFRX1TF \gr_reg[7][15]  ( .D(N831), .CK(CLK), .RN(RST_N), .Q(\GR[7][15] )
         );
  DFFRX1TF \gr_reg[7][14]  ( .D(N832), .CK(CLK), .RN(RST_N), .Q(\GR[7][14] )
         );
  DFFRX1TF \gr_reg[7][13]  ( .D(N833), .CK(CLK), .RN(RST_N), .Q(\GR[7][13] )
         );
  DFFRX1TF \gr_reg[6][15]  ( .D(N839), .CK(CLK), .RN(RST_N), .Q(\GR[6][15] )
         );
  DFFRX1TF \gr_reg[6][14]  ( .D(N840), .CK(CLK), .RN(RST_N), .Q(\GR[6][14] )
         );
  DFFRX1TF \gr_reg[6][13]  ( .D(N841), .CK(CLK), .RN(RST_N), .Q(\GR[6][13] )
         );
  DFFRX1TF \gr_reg[5][15]  ( .D(N847), .CK(CLK), .RN(RST_N), .Q(\GR[5][15] )
         );
  DFFRX1TF \gr_reg[5][14]  ( .D(N848), .CK(CLK), .RN(RST_N), .Q(\GR[5][14] )
         );
  DFFRX1TF \gr_reg[5][13]  ( .D(N849), .CK(CLK), .RN(RST_N), .Q(\GR[5][13] )
         );
  DFFRX1TF \gr_reg[4][15]  ( .D(N855), .CK(CLK), .RN(RST_N), .Q(N1389) );
  DFFRX1TF \gr_reg[4][14]  ( .D(N856), .CK(CLK), .RN(RST_N), .Q(N1390) );
  DFFRX1TF \gr_reg[4][13]  ( .D(N857), .CK(CLK), .RN(RST_N), .Q(N1391) );
  DFFRX1TF \gr_reg[3][15]  ( .D(N863), .CK(CLK), .RN(RST_N), .Q(N1386) );
  DFFRX1TF \gr_reg[3][14]  ( .D(N864), .CK(CLK), .RN(RST_N), .Q(N1387) );
  DFFRX1TF \gr_reg[3][13]  ( .D(N865), .CK(CLK), .RN(RST_N), .Q(N1388) );
  DFFRX1TF \gr_reg[2][15]  ( .D(N871), .CK(CLK), .RN(RST_N), .Q(N1383) );
  DFFRX1TF \gr_reg[2][14]  ( .D(N872), .CK(CLK), .RN(RST_N), .Q(N1384) );
  DFFRX1TF \gr_reg[2][13]  ( .D(N873), .CK(CLK), .RN(RST_N), .Q(N1385) );
  DFFRX1TF \gr_reg[1][15]  ( .D(N879), .CK(CLK), .RN(RST_N), .Q(N1375) );
  DFFRX1TF \gr_reg[1][14]  ( .D(N880), .CK(CLK), .RN(RST_N), .Q(N1376) );
  DFFRX1TF \gr_reg[1][13]  ( .D(N881), .CK(CLK), .RN(RST_N), .Q(N1377) );
  DFFRX1TF \gr_reg[0][15]  ( .D(N887), .CK(CLK), .RN(RST_N), .Q(\GR[0][15] )
         );
  DFFRX1TF \gr_reg[0][14]  ( .D(N888), .CK(CLK), .RN(RST_N), .Q(\GR[0][14] )
         );
  DFFRX1TF \gr_reg[0][13]  ( .D(N889), .CK(CLK), .RN(RST_N), .Q(\GR[0][13] )
         );
  DFFRX1TF \gr_reg[7][8]  ( .D(N838), .CK(CLK), .RN(RST_N), .Q(\GR[7][8] ) );
  DFFRX1TF \gr_reg[7][0]  ( .D(N902), .CK(CLK), .RN(RST_N), .Q(\GR[7][0] ) );
  DFFRX1TF \gr_reg[6][8]  ( .D(N846), .CK(CLK), .RN(RST_N), .Q(\GR[6][8] ) );
  DFFRX1TF \gr_reg[6][0]  ( .D(N910), .CK(CLK), .RN(RST_N), .Q(\GR[6][0] ) );
  DFFRX1TF \gr_reg[5][8]  ( .D(N854), .CK(CLK), .RN(RST_N), .Q(\GR[5][8] ) );
  DFFRX1TF \gr_reg[5][0]  ( .D(N918), .CK(CLK), .RN(RST_N), .Q(\GR[5][0] ) );
  DFFRX1TF \gr_reg[4][8]  ( .D(N862), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[8])
         );
  DFFRX1TF \gr_reg[4][0]  ( .D(N926), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[0])
         );
  DFFRX1TF \gr_reg[2][8]  ( .D(N878), .CK(CLK), .RN(RST_N), .Q(N31), .QN(N189)
         );
  DFFRX1TF \gr_reg[1][8]  ( .D(N886), .CK(CLK), .RN(RST_N), .Q(N1382) );
  DFFRX1TF \gr_reg[1][0]  ( .D(N950), .CK(CLK), .RN(RST_N), .Q(\IO_CONTROL[0] ) );
  DFFRX1TF \gr_reg[0][8]  ( .D(N894), .CK(CLK), .RN(RST_N), .Q(\GR[0][8] ) );
  DFFRX1TF \gr_reg[0][0]  ( .D(N958), .CK(CLK), .RN(RST_N), .Q(\GR[0][0] ) );
  DFFRX1TF \gr_reg[7][7]  ( .D(N895), .CK(CLK), .RN(RST_N), .Q(\GR[7][7] ) );
  DFFRX1TF \gr_reg[7][6]  ( .D(N896), .CK(CLK), .RN(RST_N), .Q(\GR[7][6] ) );
  DFFRX1TF \gr_reg[7][5]  ( .D(N897), .CK(CLK), .RN(RST_N), .Q(\GR[7][5] ) );
  DFFRX1TF \gr_reg[7][4]  ( .D(N898), .CK(CLK), .RN(RST_N), .Q(\GR[7][4] ) );
  DFFRX1TF \gr_reg[7][3]  ( .D(N899), .CK(CLK), .RN(RST_N), .Q(\GR[7][3] ) );
  DFFRX1TF \gr_reg[7][2]  ( .D(N900), .CK(CLK), .RN(RST_N), .Q(\GR[7][2] ) );
  DFFRX1TF \gr_reg[7][1]  ( .D(N901), .CK(CLK), .RN(RST_N), .Q(\GR[7][1] ) );
  DFFRX1TF \gr_reg[6][7]  ( .D(N903), .CK(CLK), .RN(RST_N), .Q(\GR[6][7] ) );
  DFFRX1TF \gr_reg[6][6]  ( .D(N904), .CK(CLK), .RN(RST_N), .Q(\GR[6][6] ) );
  DFFRX1TF \gr_reg[6][5]  ( .D(N905), .CK(CLK), .RN(RST_N), .Q(\GR[6][5] ) );
  DFFRX1TF \gr_reg[6][4]  ( .D(N906), .CK(CLK), .RN(RST_N), .Q(\GR[6][4] ) );
  DFFRX1TF \gr_reg[6][3]  ( .D(N907), .CK(CLK), .RN(RST_N), .Q(\GR[6][3] ) );
  DFFRX1TF \gr_reg[6][2]  ( .D(N908), .CK(CLK), .RN(RST_N), .Q(\GR[6][2] ) );
  DFFRX1TF \gr_reg[6][1]  ( .D(N909), .CK(CLK), .RN(RST_N), .Q(\GR[6][1] ) );
  DFFRX1TF \gr_reg[5][7]  ( .D(N911), .CK(CLK), .RN(RST_N), .Q(\GR[5][7] ) );
  DFFRX1TF \gr_reg[5][6]  ( .D(N912), .CK(CLK), .RN(RST_N), .Q(\GR[5][6] ) );
  DFFRX1TF \gr_reg[5][5]  ( .D(N913), .CK(CLK), .RN(RST_N), .Q(\GR[5][5] ) );
  DFFRX1TF \gr_reg[5][4]  ( .D(N914), .CK(CLK), .RN(RST_N), .Q(\GR[5][4] ) );
  DFFRX1TF \gr_reg[5][3]  ( .D(N915), .CK(CLK), .RN(RST_N), .Q(\GR[5][3] ) );
  DFFRX1TF \gr_reg[5][2]  ( .D(N916), .CK(CLK), .RN(RST_N), .Q(\GR[5][2] ) );
  DFFRX1TF \gr_reg[5][1]  ( .D(N917), .CK(CLK), .RN(RST_N), .Q(\GR[5][1] ) );
  DFFRX1TF \gr_reg[4][7]  ( .D(N919), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[7])
         );
  DFFRX1TF \gr_reg[4][6]  ( .D(N920), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[6])
         );
  DFFRX1TF \gr_reg[4][5]  ( .D(N921), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[5])
         );
  DFFRX1TF \gr_reg[4][4]  ( .D(N922), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[4])
         );
  DFFRX1TF \gr_reg[4][3]  ( .D(N923), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[3])
         );
  DFFRX1TF \gr_reg[4][2]  ( .D(N924), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[2])
         );
  DFFRX1TF \gr_reg[4][1]  ( .D(N925), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[1])
         );
  DFFRX1TF \gr_reg[3][7]  ( .D(N927), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[7])
         );
  DFFRX1TF \gr_reg[3][6]  ( .D(N928), .CK(CLK), .RN(RST_N), .Q(N23), .QN(N193)
         );
  DFFRX1TF \gr_reg[3][5]  ( .D(N929), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[5])
         );
  DFFRX1TF \gr_reg[3][4]  ( .D(N930), .CK(CLK), .RN(RST_N), .Q(N30), .QN(N195)
         );
  DFFRX1TF \gr_reg[3][3]  ( .D(N931), .CK(CLK), .RN(RST_N), .Q(N29), .QN(N202)
         );
  DFFRX1TF \gr_reg[2][7]  ( .D(N935), .CK(CLK), .RN(RST_N), .Q(N28), .QN(N323)
         );
  DFFRX1TF \gr_reg[2][6]  ( .D(N936), .CK(CLK), .RN(RST_N), .Q(N27), .QN(N2110) );
  DFFRX1TF \gr_reg[2][5]  ( .D(N937), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[5])
         );
  DFFRX1TF \gr_reg[2][4]  ( .D(N938), .CK(CLK), .RN(RST_N), .Q(N26), .QN(N321)
         );
  DFFRX1TF \gr_reg[2][3]  ( .D(N939), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[3])
         );
  DFFRX1TF \gr_reg[2][2]  ( .D(N940), .CK(CLK), .RN(RST_N), .Q(N25), .QN(N2170) );
  DFFRX1TF \gr_reg[2][1]  ( .D(N941), .CK(CLK), .RN(RST_N), .Q(N24), .QN(N204)
         );
  DFFRX1TF \gr_reg[1][6]  ( .D(N944), .CK(CLK), .RN(RST_N), .Q(\IO_CONTROL[6] ) );
  DFFRX1TF \gr_reg[1][5]  ( .D(N945), .CK(CLK), .RN(RST_N), .Q(\IO_CONTROL[5] ), .QN(\IO_CONTROL[5]_BAR ) );
  DFFRX1TF \gr_reg[1][1]  ( .D(N949), .CK(CLK), .RN(RST_N), .Q(\IO_CONTROL[1] ) );
  DFFRX1TF \gr_reg[0][7]  ( .D(N951), .CK(CLK), .RN(RST_N), .Q(\GR[0][7] ) );
  DFFRX1TF \gr_reg[0][6]  ( .D(N952), .CK(CLK), .RN(RST_N), .Q(\GR[0][6] ) );
  DFFRX1TF \gr_reg[0][5]  ( .D(N953), .CK(CLK), .RN(RST_N), .Q(\GR[0][5] ) );
  DFFRX1TF \gr_reg[0][4]  ( .D(N954), .CK(CLK), .RN(RST_N), .Q(\GR[0][4] ) );
  DFFRX1TF \gr_reg[0][3]  ( .D(N955), .CK(CLK), .RN(RST_N), .Q(\GR[0][3] ) );
  DFFRX1TF \gr_reg[0][2]  ( .D(N956), .CK(CLK), .RN(RST_N), .Q(\GR[0][2] ) );
  DFFRX1TF \gr_reg[0][1]  ( .D(N957), .CK(CLK), .RN(RST_N), .Q(\GR[0][1] ) );
  DFFRX2TF \gr_reg[3][9]  ( .D(N869), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[9])
         );
  DFFRX2TF \gr_reg[3][1]  ( .D(N933), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[1])
         );
  DFFRX2TF \gr_reg[3][12]  ( .D(N866), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTB[12]) );
  DFFRX2TF \gr_reg[2][0]  ( .D(N942), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[0])
         );
  DFFRX2TF \gr_reg[3][0]  ( .D(N934), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[0])
         );
  DFFRX2TF \gr_reg[3][2]  ( .D(N932), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[2])
         );
  DFFRX2TF \gr_reg[1][4]  ( .D(N946), .CK(CLK), .RN(RST_N), .Q(\IO_CONTROL[4] ) );
  DFFRX2TF \gr_reg[3][10]  ( .D(N868), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTB[10]) );
  DFFRX2TF \gr_reg[1][7]  ( .D(N943), .CK(CLK), .RN(RST_N), .Q(\IO_CONTROL[7] ) );
  DFFRX2TF \gr_reg[1][2]  ( .D(N948), .CK(CLK), .RN(RST_N), .Q(\IO_CONTROL[2] ) );
  DFFRX2TF \gr_reg[3][8]  ( .D(N870), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[8])
         );
  DFFRX2TF \gr_reg[1][3]  ( .D(N947), .CK(CLK), .RN(RST_N), .Q(\IO_CONTROL[3] ) );
  DFFRX2TF \id_ir_reg[11]  ( .D(N517), .CK(CLK), .RN(RST_N), .Q(N372), .QN(
        N560) );
  NOR2X1TF U3 ( .A(N1120), .B(N377), .Y(N606) );
  NAND2X1TF U4 ( .A(CODE_TYPE[1]), .B(N1116), .Y(N1044) );
  NAND2BX1TF U5 ( .AN(REG_A[0]), .B(REG_B[0]), .Y(SUB_X_299_4_N16) );
  NOR2X1TF U6 ( .A(N390), .B(N623), .Y(N1123) );
  CLKBUFX2TF U7 ( .A(N1041), .Y(N188) );
  CMPR32X2TF U8 ( .A(N565), .B(REG_A[15]), .C(SUB_X_299_4_N2), .CO(
        SUB_X_299_4_N1), .S(N506) );
  CLKINVX1TF U9 ( .A(N2130), .Y(N1) );
  OAI21X1TF U10 ( .A0(N804), .A1(N1), .B0(N1033), .Y(N643) );
  AOI21X1TF U11 ( .A0(REG_A[11]), .A1(N426), .B0(N771), .Y(N2) );
  NAND3X1TF U12 ( .A(N769), .B(N770), .C(N2), .Y(N1010) );
  AOI21X1TF U13 ( .A0(N614), .A1(N1091), .B0(N22), .Y(N3) );
  OAI21X1TF U14 ( .A0(N3), .A1(N1118), .B0(N607), .Y(N1040) );
  AOI21X1TF U15 ( .A0(N435), .A1(N574), .B0(N201), .Y(N4) );
  OAI2BB2XLTF U16 ( .B0(N396), .B1(N4), .A0N(N788), .A1N(N1018), .Y(N5) );
  AOI22X1TF U17 ( .A0(N616), .A1(N786), .B0(N1009), .B1(N2130), .Y(N6) );
  OAI31XLTF U18 ( .A0(N768), .A1(N407), .A2(N998), .B0(N6), .Y(N7) );
  AOI211X1TF U19 ( .A0(N604), .A1(N787), .B0(N5), .C0(N7), .Y(N8) );
  AOI22X1TF U20 ( .A0(N425), .A1(N463), .B0(N280), .B1(N497), .Y(N9) );
  AOI22X1TF U21 ( .A0(REG_A[6]), .A1(N610), .B0(N433), .B1(N396), .Y(N10) );
  AO21X1TF U22 ( .A0(N10), .A1(N615), .B0(N574), .Y(N11) );
  NAND3X1TF U23 ( .A(N8), .B(N9), .C(N11), .Y(N1080) );
  AOI2BB2X1TF U24 ( .B0(I_DATAIN[6]), .B1(N335), .A0N(N1158), .A1N(N614), .Y(
        N1700) );
  NAND4X1TF U25 ( .A(N1070), .B(N1043), .C(N1067), .D(N1063), .Y(N12) );
  NAND4BX1TF U26 ( .AN(N1072), .B(N597), .C(N601), .D(N600), .Y(N13) );
  NAND3X1TF U27 ( .A(N583), .B(N598), .C(N596), .Y(N14) );
  NOR4XLTF U28 ( .A(N1080), .B(N1058), .C(N13), .D(N14), .Y(N15) );
  NAND4X1TF U29 ( .A(N602), .B(N592), .C(N6030), .D(N15), .Y(N16) );
  NAND2X1TF U30 ( .A(N1040), .B(ZF), .Y(N17) );
  OAI31X1TF U31 ( .A0(N1053), .A1(N12), .A2(N16), .B0(N17), .Y(N287) );
  AOI21X1TF U32 ( .A0(N1125), .A1(N614), .B0(N22), .Y(N18) );
  NAND3X1TF U33 ( .A(N1124), .B(N1126), .C(N18), .Y(N223) );
  NAND3BX1TF U34 ( .AN(N91), .B(N89), .C(N90), .Y(N1166) );
  AOI2BB1X1TF U35 ( .A0N(N1024), .A1N(N804), .B0(N643), .Y(N561) );
  AOI21X1TF U36 ( .A0(REG_A[4]), .A1(N426), .B0(N971), .Y(N19) );
  NAND3X1TF U37 ( .A(N767), .B(N822), .C(N19), .Y(N1009) );
  NAND3BX1TF U38 ( .AN(N94), .B(N92), .C(N93), .Y(N1238) );
  NAND3BX1TF U39 ( .AN(N97), .B(N95), .C(N96), .Y(N1310) );
  NAND3BX1TF U40 ( .AN(N1154), .B(N545), .C(N370), .Y(N1156) );
  CLKINVX1TF U41 ( .A(N280), .Y(N20) );
  OAI22X1TF U42 ( .A0(SUB_X_299_4_N1), .A1(N20), .B0(N21), .B1(N648), .Y(N576)
         );
  CLKINVX1TF U43 ( .A(N473), .Y(N21) );
  NAND2X4TF U44 ( .A(N560), .B(CODE_TYPE[2]), .Y(N1091) );
  OR3X2TF U45 ( .A(REG_B[3]), .B(REG_B[2]), .C(N1014), .Y(N608) );
  AOI21X2TF U46 ( .A0(N578), .A1(REG_B[0]), .B0(N577), .Y(N601) );
  AOI22XLTF U47 ( .A0(N292), .A1(\IO_CONTROL[2] ), .B0(N270), .B1(
        IO_DATAOUTB[2]), .Y(N1176) );
  AOI22XLTF U48 ( .A0(N310), .A1(\IO_CONTROL[2] ), .B0(N268), .B1(
        IO_DATAOUTB[2]), .Y(N1248) );
  AOI22XLTF U49 ( .A0(N313), .A1(\IO_CONTROL[2] ), .B0(N273), .B1(
        IO_DATAOUTB[2]), .Y(N1320) );
  INVX1TF U59 ( .A(N561), .Y(N541) );
  OA21XLTF U60 ( .A0(N1119), .A1(N1128), .B0(N1150), .Y(N1152) );
  OAI21XLTF U61 ( .A0(N736), .A1(I_ADDR[6]), .B0(N739), .Y(N737) );
  NAND2X1TF U62 ( .A(N584), .B(N1042), .Y(N594) );
  OAI2BB1X1TF U63 ( .A0N(N612), .A1N(N606), .B0(N437), .Y(N1032) );
  NOR2X1TF U64 ( .A(N453), .B(N424), .Y(N1084) );
  OR2X2TF U65 ( .A(N665), .B(N1044), .Y(N1033) );
  NAND2XLTF U66 ( .A(REG_A[10]), .B(N2220), .Y(N635) );
  NAND2X1TF U67 ( .A(REG_A[11]), .B(N2220), .Y(N639) );
  OAI21XLTF U68 ( .A0(I_ADDR[1]), .A1(I_ADDR[2]), .B0(N727), .Y(N725) );
  OR3X1TF U69 ( .A(N91), .B(N89), .C(N90), .Y(N1159) );
  OR3X1TF U70 ( .A(N97), .B(N95), .C(N404), .Y(N1304) );
  OR3X1TF U71 ( .A(N94), .B(N92), .C(N403), .Y(N1232) );
  OR3X1TF U72 ( .A(N89), .B(N90), .C(N374), .Y(N1162) );
  AOI21X2TF U73 ( .A0(N504), .A1(N280), .B0(N4570), .Y(N6030) );
  AOI211X1TF U74 ( .A0(N346), .A1(D_ADDR[3]), .B0(N729), .C0(N728), .Y(N721)
         );
  AOI211X1TF U75 ( .A0(N346), .A1(D_ADDR[5]), .B0(N735), .C0(N734), .Y(N719)
         );
  AOI211X1TF U76 ( .A0(N346), .A1(D_ADDR[7]), .B0(N741), .C0(N740), .Y(N717)
         );
  AOI21X1TF U77 ( .A0(D_ADDR[8]), .A1(N346), .B0(N747), .Y(N713) );
  AOI21X1TF U78 ( .A0(D_ADDR[2]), .A1(N346), .B0(N726), .Y(N722) );
  AOI211X1TF U79 ( .A0(N346), .A1(D_ADDR[9]), .B0(N657), .C0(N656), .Y(N775)
         );
  AOI21X1TF U80 ( .A0(D_ADDR[6]), .A1(N346), .B0(N738), .Y(N718) );
  AOI21X1TF U81 ( .A0(D_ADDR[4]), .A1(N346), .B0(N732), .Y(N720) );
  OR2X2TF U82 ( .A(N680), .B(N703), .Y(N677) );
  OR2X2TF U83 ( .A(N678), .B(N703), .Y(N676) );
  OR2X2TF U84 ( .A(N700), .B(N707), .Y(N701) );
  OR2X2TF U85 ( .A(N697), .B(N678), .Y(N671) );
  OR2X2TF U86 ( .A(N680), .B(N700), .Y(N675) );
  OR2X2TF U87 ( .A(N678), .B(N708), .Y(N679) );
  OR2X2TF U88 ( .A(N708), .B(N705), .Y(N706) );
  OR2X2TF U89 ( .A(N703), .B(N707), .Y(N704) );
  OR2X2TF U90 ( .A(N697), .B(N707), .Y(N698) );
  OR2X2TF U91 ( .A(N697), .B(N705), .Y(N695) );
  OR2X2TF U92 ( .A(N700), .B(N705), .Y(N699) );
  OR2X2TF U93 ( .A(N680), .B(N708), .Y(N689) );
  AOI22X1TF U94 ( .A0(N326), .A1(N175), .B0(N347), .B1(N212), .Y(N1107) );
  AOI22X1TF U95 ( .A0(N325), .A1(N185), .B0(N1112), .B1(N222), .Y(N1097) );
  AOI22X1TF U96 ( .A0(N326), .A1(N174), .B0(N1112), .B1(N211), .Y(N1108) );
  AOI22X1TF U97 ( .A0(N325), .A1(N180), .B0(N1112), .B1(N217), .Y(N1102) );
  AOI22X1TF U98 ( .A0(N325), .A1(N173), .B0(N1112), .B1(N210), .Y(N1109) );
  AOI22X1TF U99 ( .A0(N326), .A1(N179), .B0(N347), .B1(N216), .Y(N1103) );
  AOI22X1TF U100 ( .A0(N325), .A1(N171), .B0(N1112), .B1(N208), .Y(N1111) );
  AOI22X1TF U101 ( .A0(N326), .A1(N182), .B0(N1112), .B1(N219), .Y(N1100) );
  AOI22X1TF U102 ( .A0(N326), .A1(N183), .B0(N347), .B1(N220), .Y(N1099) );
  AOI22X1TF U103 ( .A0(N325), .A1(N172), .B0(N1112), .B1(N209), .Y(N1110) );
  AOI22X1TF U104 ( .A0(N326), .A1(N177), .B0(N347), .B1(N214), .Y(N1105) );
  AOI22X1TF U105 ( .A0(N325), .A1(N184), .B0(N1112), .B1(N221), .Y(N1098) );
  AOI22X1TF U106 ( .A0(N326), .A1(N178), .B0(N347), .B1(N215), .Y(N1104) );
  AOI22X1TF U107 ( .A0(N325), .A1(N176), .B0(N1112), .B1(N213), .Y(N1106) );
  OAI21XLTF U108 ( .A0(N406), .A1(N234), .B0(N1131), .Y(N486) );
  AOI22X1TF U109 ( .A0(N326), .A1(N181), .B0(N347), .B1(N218), .Y(N1101) );
  AOI22X1TF U110 ( .A0(N325), .A1(N170), .B0(N1112), .B1(N207), .Y(N1113) );
  INVX1TF U111 ( .A(N693), .Y(N692) );
  NAND4XLTF U112 ( .A(N647), .B(N646), .C(N648), .D(N373), .Y(N575) );
  INVX2TF U113 ( .A(N1084), .Y(N198) );
  OAI211X1TF U114 ( .A0(N1128), .A1(N1094), .B0(N1095), .C0(N1096), .Y(N1114)
         );
  NAND3XLTF U115 ( .A(N760), .B(N759), .C(N1153), .Y(NEXT_STATE[2]) );
  CLKINVX2TF U116 ( .A(N1031), .Y(N1035) );
  INVX2TF U117 ( .A(N1033), .Y(N200) );
  NAND2XLTF U118 ( .A(REG_B[3]), .B(N790), .Y(N791) );
  OR2X2TF U119 ( .A(N690), .B(N654), .Y(N345) );
  OAI31XLTF U120 ( .A0(STATE[3]), .A1(INSTR_OVER), .A2(N758), .B0(N757), .Y(
        N760) );
  NOR2X4TF U121 ( .A(N662), .B(N1127), .Y(N694) );
  AOI22X1TF U122 ( .A0(N316), .A1(\GR[0][2] ), .B0(N274), .B1(N25), .Y(N1247)
         );
  AOI22X1TF U123 ( .A0(N314), .A1(\GR[0][2] ), .B0(N276), .B1(N25), .Y(N1319)
         );
  AOI22X1TF U124 ( .A0(N231), .A1(IO_OFFSET[6]), .B0(N281), .B1(\GR[6][6] ), 
        .Y(N1193) );
  AOI22X1TF U125 ( .A0(N231), .A1(IO_OFFSET[5]), .B0(N281), .B1(\GR[6][5] ), 
        .Y(N1189) );
  AOI22X1TF U126 ( .A0(N229), .A1(\GR[0][6] ), .B0(N283), .B1(N27), .Y(N1191)
         );
  AND2X2TF U127 ( .A(N1093), .B(N1042), .Y(N609) );
  AOI22X1TF U128 ( .A0(N1234), .A1(N1389), .B0(N285), .B1(\GR[6][15] ), .Y(
        N1301) );
  OAI21XLTF U129 ( .A0(N730), .A1(I_ADDR[4]), .B0(N733), .Y(N731) );
  AOI22X1TF U130 ( .A0(N1234), .A1(IO_OFFSET[1]), .B0(N285), .B1(\GR[6][1] ), 
        .Y(N1245) );
  AOI22X1TF U131 ( .A0(N229), .A1(\GR[0][5] ), .B0(N283), .B1(IO_DATAOUTA[5]), 
        .Y(N1187) );
  AOI22X1TF U132 ( .A0(N1234), .A1(IO_OFFSET[9]), .B0(N285), .B1(\GR[6][9] ), 
        .Y(N1277) );
  AOI22X1TF U133 ( .A0(N1234), .A1(IO_OFFSET[5]), .B0(N285), .B1(\GR[6][5] ), 
        .Y(N1261) );
  AOI22X1TF U134 ( .A0(N1234), .A1(N1390), .B0(N285), .B1(\GR[6][14] ), .Y(
        N1297) );
  AOI22X1TF U135 ( .A0(N229), .A1(\GR[0][2] ), .B0(N283), .B1(N25), .Y(N1175)
         );
  AOI22X1TF U136 ( .A0(N1306), .A1(IO_OFFSET[8]), .B0(N290), .B1(\GR[6][8] ), 
        .Y(N1345) );
  AOI22X1TF U137 ( .A0(N229), .A1(\GR[0][12] ), .B0(N283), .B1(N34), .Y(N1215)
         );
  AOI22X1TF U138 ( .A0(N1306), .A1(IO_OFFSET[9]), .B0(N290), .B1(\GR[6][9] ), 
        .Y(N1349) );
  AOI22X1TF U139 ( .A0(N231), .A1(IO_OFFSET[2]), .B0(N281), .B1(\GR[6][2] ), 
        .Y(N1177) );
  AOI22X1TF U140 ( .A0(N1306), .A1(N1394), .B0(N290), .B1(\GR[6][10] ), .Y(
        N1353) );
  AOI22X1TF U141 ( .A0(N231), .A1(N1392), .B0(N281), .B1(\GR[6][12] ), .Y(
        N1217) );
  AOI22X1TF U142 ( .A0(N229), .A1(\GR[0][1] ), .B0(N283), .B1(N24), .Y(N1171)
         );
  AOI22X1TF U143 ( .A0(N1306), .A1(N1392), .B0(N290), .B1(\GR[6][12] ), .Y(
        N1361) );
  AOI22X1TF U144 ( .A0(N1306), .A1(N1390), .B0(N290), .B1(\GR[6][14] ), .Y(
        N1369) );
  AOI22X1TF U145 ( .A0(N231), .A1(IO_OFFSET[1]), .B0(N281), .B1(\GR[6][1] ), 
        .Y(N1173) );
  AOI22X1TF U146 ( .A0(N1306), .A1(N1391), .B0(N290), .B1(\GR[6][13] ), .Y(
        N1365) );
  AOI22X1TF U147 ( .A0(N231), .A1(IO_OFFSET[0]), .B0(N281), .B1(\GR[6][0] ), 
        .Y(N1169) );
  AOI22X1TF U148 ( .A0(N1234), .A1(IO_OFFSET[0]), .B0(N285), .B1(\GR[6][0] ), 
        .Y(N1241) );
  AOI22X1TF U149 ( .A0(N229), .A1(\GR[0][0] ), .B0(N283), .B1(IO_DATAOUTA[0]), 
        .Y(N1167) );
  OR2X1TF U150 ( .A(N761), .B(N1124), .Y(NEXT_STATE[3]) );
  OR3X1TF U151 ( .A(N409), .B(N370), .C(N1154), .Y(N1153) );
  INVX2TF U152 ( .A(REG_B[2]), .Y(N197) );
  INVX2TF U153 ( .A(N384), .Y(N2100) );
  OR3X1TF U154 ( .A(N91), .B(N89), .C(N380), .Y(N1160) );
  OR3X1TF U155 ( .A(N91), .B(N90), .C(N381), .Y(N1161) );
  OR3X1TF U156 ( .A(N89), .B(N374), .C(N380), .Y(N1163) );
  OR3X1TF U157 ( .A(N94), .B(N92), .C(N93), .Y(N1231) );
  NOR2X4TF U158 ( .A(N406), .B(N371), .Y(N807) );
  OR3X1TF U159 ( .A(N94), .B(N93), .C(N382), .Y(N1233) );
  OR3X1TF U160 ( .A(N92), .B(N376), .C(N403), .Y(N1235) );
  OR3X1TF U161 ( .A(N95), .B(N375), .C(N404), .Y(N1307) );
  OR3X1TF U162 ( .A(N97), .B(N95), .C(N96), .Y(N1303) );
  OR3X1TF U163 ( .A(N97), .B(N96), .C(N383), .Y(N1305) );
  INVX2TF U164 ( .A(N189), .Y(IO_DATAOUTA[8]) );
  INVX2TF U165 ( .A(N191), .Y(IO_DATAOUTA[10]) );
  INVX2TF U166 ( .A(N193), .Y(IO_DATAOUTB[6]) );
  INVX2TF U167 ( .A(N195), .Y(IO_DATAOUTB[4]) );
  INVX2TF U168 ( .A(N1084), .Y(N199) );
  INVX2TF U169 ( .A(N1033), .Y(N201) );
  INVX2TF U170 ( .A(N202), .Y(IO_DATAOUTB[3]) );
  INVX2TF U171 ( .A(N204), .Y(IO_DATAOUTA[1]) );
  INVX2TF U172 ( .A(N206), .Y(IO_DATAOUTA[12]) );
  INVX2TF U173 ( .A(N2080), .Y(IO_DATAOUTB[11]) );
  INVX2TF U174 ( .A(N2110), .Y(IO_DATAOUTA[6]) );
  INVX2TF U175 ( .A(N608), .Y(N2130) );
  INVX2TF U176 ( .A(N608), .Y(N2140) );
  INVX2TF U177 ( .A(N594), .Y(N2150) );
  INVX2TF U178 ( .A(N594), .Y(N2160) );
  INVX2TF U179 ( .A(N2170), .Y(IO_DATAOUTA[2]) );
  INVX2TF U180 ( .A(N1153), .Y(N2190) );
  INVX2TF U181 ( .A(N1153), .Y(N2200) );
  INVX2TF U182 ( .A(N804), .Y(N2210) );
  INVX2TF U183 ( .A(N804), .Y(N2220) );
  INVX2TF U184 ( .A(N223), .Y(N224) );
  INVX2TF U185 ( .A(N223), .Y(N225) );
  INVX2TF U186 ( .A(N1114), .Y(N226) );
  INVX2TF U187 ( .A(N226), .Y(N227) );
  INVX2TF U188 ( .A(N226), .Y(N228) );
  INVX2TF U189 ( .A(N1159), .Y(N229) );
  INVX2TF U190 ( .A(N1159), .Y(N230) );
  INVX2TF U191 ( .A(N1162), .Y(N231) );
  INVX2TF U192 ( .A(N1162), .Y(N232) );
  INVX2TF U193 ( .A(N1152), .Y(N233) );
  INVX2TF U194 ( .A(N1152), .Y(N234) );
  INVX2TF U195 ( .A(N706), .Y(N235) );
  INVX2TF U196 ( .A(N706), .Y(N236) );
  INVX2TF U197 ( .A(N695), .Y(N237) );
  INVX2TF U198 ( .A(N695), .Y(N238) );
  INVX2TF U199 ( .A(N689), .Y(N239) );
  INVX2TF U200 ( .A(N689), .Y(N240) );
  INVX2TF U201 ( .A(N679), .Y(N241) );
  INVX2TF U202 ( .A(N679), .Y(N242) );
  INVX2TF U203 ( .A(N676), .Y(N243) );
  INVX2TF U204 ( .A(N676), .Y(N244) );
  INVX2TF U205 ( .A(N671), .Y(N245) );
  INVX2TF U206 ( .A(N671), .Y(N246) );
  INVX2TF U207 ( .A(N677), .Y(N2470) );
  INVX2TF U208 ( .A(N677), .Y(N2480) );
  INVX2TF U209 ( .A(N701), .Y(N2490) );
  INVX2TF U210 ( .A(N701), .Y(N2500) );
  INVX2TF U211 ( .A(N704), .Y(N2510) );
  INVX2TF U212 ( .A(N704), .Y(N2520) );
  INVX2TF U213 ( .A(N698), .Y(N2530) );
  INVX2TF U214 ( .A(N698), .Y(N263) );
  INVX2TF U215 ( .A(N699), .Y(N264) );
  INVX2TF U216 ( .A(N699), .Y(N265) );
  INVX2TF U217 ( .A(N675), .Y(N266) );
  INVX2TF U218 ( .A(N675), .Y(N267) );
  INVX2TF U219 ( .A(N1238), .Y(N268) );
  INVX2TF U220 ( .A(N1238), .Y(N269) );
  INVX2TF U221 ( .A(N1166), .Y(N270) );
  INVX2TF U222 ( .A(N1166), .Y(N271) );
  INVX2TF U223 ( .A(N1310), .Y(N272) );
  INVX2TF U224 ( .A(N1310), .Y(N273) );
  INVX2TF U225 ( .A(N1232), .Y(N274) );
  INVX2TF U226 ( .A(N1232), .Y(N275) );
  INVX2TF U227 ( .A(N1304), .Y(N276) );
  INVX2TF U228 ( .A(N1304), .Y(N277) );
  INVX2TF U229 ( .A(N1032), .Y(N278) );
  INVX2TF U230 ( .A(N278), .Y(N279) );
  INVX2TF U231 ( .A(N278), .Y(N280) );
  AOI22XLTF U232 ( .A0(N1026), .A1(N987), .B0(N1031), .B1(N986), .Y(N540) );
  NOR2X2TF U233 ( .A(N614), .B(N384), .Y(N1122) );
  OAI31X4TF U234 ( .A0(N1129), .A1(N1128), .A2(N1127), .B0(N1140), .Y(N1133)
         );
  OAI21X1TF U235 ( .A0(N545), .A1(N754), .B0(N645), .Y(N165) );
  INVX2TF U236 ( .A(N1163), .Y(N281) );
  INVX2TF U237 ( .A(N1163), .Y(N282) );
  INVX2TF U238 ( .A(N1160), .Y(N283) );
  INVX2TF U239 ( .A(N1160), .Y(N284) );
  INVX2TF U240 ( .A(N1235), .Y(N285) );
  INVX2TF U241 ( .A(N1235), .Y(N286) );
  INVX2TF U242 ( .A(N1307), .Y(N290) );
  INVX2TF U243 ( .A(N1307), .Y(N291) );
  INVX2TF U244 ( .A(N1161), .Y(N292) );
  INVX2TF U245 ( .A(N1161), .Y(N309) );
  INVX2TF U246 ( .A(N1233), .Y(N310) );
  INVX2TF U247 ( .A(N1233), .Y(N311) );
  INVX2TF U248 ( .A(N1305), .Y(N312) );
  INVX2TF U249 ( .A(N1305), .Y(N313) );
  INVX2TF U250 ( .A(N1303), .Y(N314) );
  INVX2TF U251 ( .A(N1303), .Y(N315) );
  INVX2TF U252 ( .A(N1231), .Y(N316) );
  INVX2TF U253 ( .A(N1231), .Y(N317) );
  NAND2X2TF U254 ( .A(N757), .B(N752), .Y(N690) );
  NOR3X2TF U255 ( .A(N545), .B(N546), .C(STATE[1]), .Y(N757) );
  INVX2TF U256 ( .A(N188), .Y(N319) );
  INVX2TF U257 ( .A(N188), .Y(N320) );
  INVX2TF U258 ( .A(N321), .Y(IO_DATAOUTA[4]) );
  INVX2TF U259 ( .A(N323), .Y(IO_DATAOUTA[7]) );
  INVX2TF U260 ( .A(N1095), .Y(N325) );
  INVX2TF U261 ( .A(N1095), .Y(N326) );
  INVX2TF U262 ( .A(N327), .Y(IO_DATAOUTA[9]) );
  INVXLTF U263 ( .A(N1024), .Y(N330) );
  INVX2TF U264 ( .A(N1024), .Y(N616) );
  NAND3X1TF U265 ( .A(N407), .B(N197), .C(N790), .Y(N1024) );
  INVX2TF U266 ( .A(N1081), .Y(N331) );
  OAI21X1TF U267 ( .A0(N591), .A1(N331), .B0(N590), .Y(N318) );
  OA22X1TF U268 ( .A0(N601), .A1(N1078), .B0(N1070), .B1(N198), .Y(N1045) );
  NAND2X1TF U269 ( .A(N611), .B(N607), .Y(N1078) );
  INVX2TF U270 ( .A(N807), .Y(N332) );
  INVX2TF U271 ( .A(N807), .Y(N993) );
  INVX2TF U272 ( .A(N968), .Y(N333) );
  CLKBUFX2TF U273 ( .A(N593), .Y(N334) );
  NOR2BX1TF U274 ( .AN(N584), .B(N1125), .Y(N593) );
  INVX2TF U275 ( .A(N1156), .Y(N335) );
  CLKBUFX2TF U276 ( .A(N724), .Y(N336) );
  NOR2X2TF U277 ( .A(N708), .B(N707), .Y(N724) );
  CLKBUFX2TF U278 ( .A(N702), .Y(N337) );
  NOR2X2TF U279 ( .A(N703), .B(N705), .Y(N702) );
  CLKBUFX2TF U280 ( .A(N673), .Y(N339) );
  NOR2X2TF U281 ( .A(N697), .B(N680), .Y(N673) );
  CLKBUFX2TF U282 ( .A(N674), .Y(N340) );
  NOR2X2TF U283 ( .A(N678), .B(N700), .Y(N674) );
  CLKBUFX2TF U284 ( .A(N431), .Y(N341) );
  CLKBUFX2TF U285 ( .A(N1308), .Y(N431) );
  CLKBUFX2TF U286 ( .A(N429), .Y(N342) );
  CLKBUFX2TF U287 ( .A(N1236), .Y(N429) );
  INVX2TF U288 ( .A(N969), .Y(N343) );
  CLKBUFX2TF U289 ( .A(N990), .Y(N426) );
  NOR3BXLTF U290 ( .AN(INSTR_OVER), .B(N758), .C(N690), .Y(N167) );
  OAI21XLTF U291 ( .A0(N758), .A1(N751), .B0(N750), .Y(NEXT_STATE[0]) );
  AOI22XLTF U292 ( .A0(N496), .A1(N279), .B0(N462), .B1(N580), .Y(N581) );
  AOI22XLTF U293 ( .A0(N2140), .A1(N963), .B0(N461), .B1(N580), .Y(N533) );
  AOI21XLTF U294 ( .A0(N468), .A1(N580), .B0(N512), .Y(N514) );
  INVX2TF U295 ( .A(N983), .Y(N344) );
  NOR2BX2TF U296 ( .AN(N22), .B(CODE_TYPE[3]), .Y(N612) );
  INVX2TF U297 ( .A(N345), .Y(N346) );
  AOI21XLTF U298 ( .A0(D_ADDR[1]), .A1(N346), .B0(N655), .Y(N776) );
  NOR2X2TF U299 ( .A(N197), .B(REG_B[3]), .Y(N988) );
  INVX2TF U300 ( .A(N1096), .Y(N347) );
  AOI32X1TF U301 ( .A0(N1115), .A1(N1124), .A2(N1093), .B0(N1092), .B1(N1124), 
        .Y(N1096) );
  NAND3X2TF U302 ( .A(N606), .B(N1093), .C(N1124), .Y(N1041) );
  CLKBUFX2TF U303 ( .A(N1164), .Y(N349) );
  CLKBUFX2TF U304 ( .A(N1306), .Y(N350) );
  CLKBUFX2TF U305 ( .A(N1234), .Y(N351) );
  NOR4X4TF U306 ( .A(N370), .B(N395), .C(N545), .D(STATE[3]), .Y(N1124) );
  XOR2X1TF U307 ( .A(REG_A[0]), .B(REG_B[0]), .Y(N491) );
  CMPR32X2TF U308 ( .A(N352), .B(REG_A[3]), .C(SUB_X_299_4_N14), .CO(
        SUB_X_299_4_N13), .S(N494) );
  ADDFHX2TF U309 ( .A(N571), .B(REG_A[9]), .CI(SUB_X_299_4_N8), .CO(
        SUB_X_299_4_N7), .S(N500) );
  ADDFHX2TF U310 ( .A(N5760), .B(REG_A[4]), .CI(SUB_X_299_4_N13), .CO(
        SUB_X_299_4_N12), .S(N495) );
  XOR2X4TF U311 ( .A(N592), .B(N586), .Y(N591) );
  CLKXOR2X2TF U312 ( .A(N6030), .B(N585), .Y(N586) );
  OR2X2TF U313 ( .A(N451), .B(CODE_TYPE[3]), .Y(N663) );
  NAND2X1TF U314 ( .A(N406), .B(REG_B[0]), .Y(N968) );
  NAND2X2TF U315 ( .A(N472), .B(N425), .Y(N550) );
  NAND3X1TF U316 ( .A(N441), .B(N440), .C(N648), .Y(N580) );
  NAND2X1TF U317 ( .A(N372), .B(CODE_TYPE[1]), .Y(N623) );
  OAI22X1TF U318 ( .A0(ZF), .A1(N662), .B0(CF), .B1(N1091), .Y(N649) );
  INVX2TF U319 ( .A(N1015), .Y(N615) );
  AOI21X4TF U320 ( .A0(N506), .A1(N280), .B0(N552), .Y(N592) );
  INVX2TF U321 ( .A(N983), .Y(N610) );
  NAND2X1TF U322 ( .A(N696), .B(N381), .Y(N705) );
  NAND2X1TF U323 ( .A(N89), .B(N696), .Y(N707) );
  NAND2X1TF U324 ( .A(N381), .B(N672), .Y(N678) );
  NAND2X1TF U325 ( .A(N89), .B(N672), .Y(N680) );
  INVX2TF U326 ( .A(N694), .Y(N691) );
  NAND2X1TF U327 ( .A(N560), .B(N1115), .Y(N662) );
  NOR2X1TF U328 ( .A(N424), .B(N1088), .Y(N584) );
  OAI21X2TF U329 ( .A0(N1087), .A1(N1094), .B0(N647), .Y(N1015) );
  INVX2TF U330 ( .A(N1093), .Y(N1127) );
  NOR2X1TF U331 ( .A(CODE_TYPE[2]), .B(N377), .Y(N1115) );
  NOR2X1TF U332 ( .A(N1116), .B(N1115), .Y(N1129) );
  NOR3X1TF U333 ( .A(N759), .B(N975), .C(N1127), .Y(N603) );
  AOI21X1TF U334 ( .A0(N691), .A1(N693), .B0(N690), .Y(N696) );
  OAI22X1TF U335 ( .A0(N690), .A1(N693), .B0(N691), .B1(N668), .Y(N672) );
  AOI21X2TF U336 ( .A0(N505), .A1(N280), .B0(N4640), .Y(N602) );
  CLKBUFX2TF U337 ( .A(N1079), .Y(N424) );
  OR2X2TF U338 ( .A(N759), .B(N409), .Y(N1079) );
  CLKBUFX2TF U339 ( .A(N580), .Y(N425) );
  NOR2X2TF U340 ( .A(CODE_TYPE[3]), .B(N2100), .Y(N1093) );
  NOR2X2TF U341 ( .A(CODE_TYPE[1]), .B(N1091), .Y(N1042) );
  INVX2TF U342 ( .A(N1096), .Y(N1112) );
  NAND2X1TF U343 ( .A(N90), .B(N91), .Y(N708) );
  NAND2X1TF U344 ( .A(N90), .B(N374), .Y(N700) );
  NAND2X1TF U345 ( .A(N380), .B(N374), .Y(N697) );
  INVX2TF U346 ( .A(N690), .Y(N670) );
  NAND2X1TF U347 ( .A(N91), .B(N380), .Y(N703) );
  NAND2X1TF U348 ( .A(STATE[3]), .B(N757), .Y(N668) );
  INVX2TF U349 ( .A(N424), .Y(N607) );
  NAND2X1TF U350 ( .A(N372), .B(N390), .Y(N1120) );
  AOI211XLTF U351 ( .A0(N22), .A1(N1123), .B0(CODE_TYPE[3]), .C0(N1117), .Y(
        N1119) );
  AOI221XLTF U352 ( .A0(N560), .A1(N416), .B0(N372), .B1(NF), .C0(CODE_TYPE[1]), .Y(N650) );
  INVX2TF U353 ( .A(N1156), .Y(N1158) );
  NAND2X1TF U354 ( .A(N752), .B(STATE[1]), .Y(N1154) );
  INVX2TF U355 ( .A(N668), .Y(N669) );
  NAND3X1TF U356 ( .A(STATE[3]), .B(STATE[1]), .C(N370), .Y(N759) );
  NOR2X1TF U357 ( .A(N1125), .B(N1127), .Y(N611) );
  NAND3X1TF U358 ( .A(CODE_TYPE[2]), .B(N377), .C(N372), .Y(N1125) );
  AO22X1TF U359 ( .A0(N600), .A1(CF_BUF), .B0(N1040), .B1(CF), .Y(N289) );
  AO22X1TF U360 ( .A0(N319), .A1(N175), .B0(N1041), .B1(SMDR[10]), .Y(N303) );
  AO22X1TF U361 ( .A0(N319), .A1(N174), .B0(N1041), .B1(SMDR[11]), .Y(N304) );
  AO22X1TF U362 ( .A0(N319), .A1(N177), .B0(N1041), .B1(SMDR[8]), .Y(N301) );
  AO22X1TF U363 ( .A0(N319), .A1(N178), .B0(N1041), .B1(SMDR[7]), .Y(N300) );
  AO22X1TF U364 ( .A0(N319), .A1(N180), .B0(N1041), .B1(SMDR[5]), .Y(N298) );
  AO22X1TF U365 ( .A0(N319), .A1(N176), .B0(N1041), .B1(SMDR[9]), .Y(N302) );
  AO22X1TF U366 ( .A0(N319), .A1(N184), .B0(N1041), .B1(SMDR[1]), .Y(N294) );
  AO22X1TF U367 ( .A0(N319), .A1(N173), .B0(N1041), .B1(SMDR[12]), .Y(N305) );
  AO22X1TF U368 ( .A0(N320), .A1(N172), .B0(N188), .B1(SMDR[13]), .Y(N306) );
  AO22X1TF U369 ( .A0(N320), .A1(N182), .B0(N188), .B1(SMDR[3]), .Y(N296) );
  AO22X1TF U370 ( .A0(N320), .A1(N171), .B0(N188), .B1(SMDR[14]), .Y(N307) );
  AO22X1TF U371 ( .A0(N320), .A1(N170), .B0(N188), .B1(SMDR[15]), .Y(N308) );
  AO22X1TF U372 ( .A0(N320), .A1(N179), .B0(N188), .B1(SMDR[6]), .Y(N299) );
  AO22X1TF U373 ( .A0(N320), .A1(N185), .B0(N188), .B1(SMDR[0]), .Y(N293) );
  AO22X1TF U374 ( .A0(N320), .A1(N181), .B0(N188), .B1(SMDR[4]), .Y(N297) );
  AO22X1TF U375 ( .A0(N320), .A1(N183), .B0(N188), .B1(SMDR[2]), .Y(N295) );
  NOR3X1TF U376 ( .A(CODE_TYPE[1]), .B(N1120), .C(N1127), .Y(N758) );
  AOI22XLTF U377 ( .A0(N312), .A1(\IO_CONTROL[5] ), .B0(N272), .B1(
        IO_DATAOUTB[5]), .Y(N1332) );
  AOI22XLTF U378 ( .A0(N312), .A1(\IO_CONTROL[6] ), .B0(N272), .B1(N23), .Y(
        N1336) );
  AOI22XLTF U379 ( .A0(N310), .A1(\IO_CONTROL[5] ), .B0(N268), .B1(
        IO_DATAOUTB[5]), .Y(N1260) );
  AOI22XLTF U380 ( .A0(N292), .A1(\IO_CONTROL[5] ), .B0(N270), .B1(
        IO_DATAOUTB[5]), .Y(N1188) );
  AOI22XLTF U381 ( .A0(N310), .A1(\IO_CONTROL[6] ), .B0(N268), .B1(N23), .Y(
        N1264) );
  AOI22XLTF U382 ( .A0(N292), .A1(\IO_CONTROL[6] ), .B0(N270), .B1(N23), .Y(
        N1192) );
  OAI2BB2XLTF U383 ( .B0(N370), .B1(N1154), .A0N(N545), .A1N(N756), .Y(
        NEXT_STATE[1]) );
  AOI2BB2X1TF U384 ( .B0(N225), .B1(N259), .A0N(N407), .A1N(N233), .Y(N1134)
         );
  NAND2X1TF U385 ( .A(N1118), .B(N1124), .Y(N1150) );
  NOR2X1TF U386 ( .A(N1120), .B(N614), .Y(N1121) );
  OAI2BB2XLTF U387 ( .B0(N2190), .B1(N383), .A0N(N2200), .A1N(I_DATAIN[0]), 
        .Y(N508) );
  OAI2BB2XLTF U388 ( .B0(N2190), .B1(N404), .A0N(N2200), .A1N(I_DATAIN[1]), 
        .Y(N507) );
  OAI2BB2XLTF U389 ( .B0(N2190), .B1(N375), .A0N(N2200), .A1N(I_DATAIN[2]), 
        .Y(N5060) );
  OAI2BB2XLTF U390 ( .B0(N2190), .B1(N382), .A0N(N2200), .A1N(I_DATAIN[4]), 
        .Y(N5040) );
  OAI2BB2XLTF U391 ( .B0(N2190), .B1(N376), .A0N(N2200), .A1N(I_DATAIN[6]), 
        .Y(N5020) );
  OAI2BB2XLTF U392 ( .B0(N2200), .B1(N403), .A0N(N2200), .A1N(I_DATAIN[5]), 
        .Y(N5030) );
  OAI2BB2XLTF U393 ( .B0(N1158), .B1(N380), .A0N(N1158), .A1N(I_DATAIN[1]), 
        .Y(N519) );
  OAI2BB2XLTF U394 ( .B0(N1158), .B1(N377), .A0N(N1158), .A1N(I_DATAIN[4]), 
        .Y(N516) );
  OAI2BB2XLTF U395 ( .B0(N1158), .B1(N381), .A0N(N1158), .A1N(I_DATAIN[0]), 
        .Y(N520) );
  OAI2BB2XLTF U396 ( .B0(N1158), .B1(N374), .A0N(N1158), .A1N(I_DATAIN[2]), 
        .Y(N518) );
  OAI2BB2XLTF U397 ( .B0(N1158), .B1(N390), .A0N(N335), .A1N(I_DATAIN[5]), .Y(
        N515) );
  AOI22XLTF U398 ( .A0(IS_I_ADDR), .A1(N1128), .B0(N749), .B1(N370), .Y(N661)
         );
  AO21X1TF U399 ( .A0(N660), .A1(N659), .B0(N748), .Y(N960) );
  AOI2BB2X2TF U400 ( .B0(D_DATAIN[1]), .B1(N694), .A0N(N2620), .A1N(N693), .Y(
        N710) );
  AOI2BB2X2TF U401 ( .B0(D_DATAIN[4]), .B1(N694), .A0N(N2610), .A1N(N693), .Y(
        N714) );
  AOI2BB2X2TF U402 ( .B0(D_DATAIN[2]), .B1(N694), .A0N(N2580), .A1N(N693), .Y(
        N711) );
  AOI2BB2X2TF U403 ( .B0(D_DATAIN[6]), .B1(N694), .A0N(N2570), .A1N(N693), .Y(
        N716) );
  AOI2BB2X2TF U405 ( .B0(D_DATAIN[5]), .B1(N694), .A0N(N2600), .A1N(N693), .Y(
        N715) );
  AOI2BB2X2TF U406 ( .B0(D_DATAIN[3]), .B1(N694), .A0N(N2590), .A1N(N693), .Y(
        N712) );
  AOI2BB2X2TF U407 ( .B0(D_DATAIN[7]), .B1(N694), .A0N(N2560), .A1N(N693), .Y(
        N723) );
  AO21X1TF U408 ( .A0(N1075), .A1(N1072), .B0(N1071), .Y(N418) );
  NAND2X2TF U409 ( .A(N406), .B(N371), .Y(N804) );
  OAI21X1TF U410 ( .A0(N619), .A1(N1116), .B0(N22), .Y(N439) );
  NOR2X1TF U411 ( .A(N344), .B(N280), .Y(N646) );
  AOI211X1TF U412 ( .A0(START), .A1(N749), .B0(N761), .C0(N748), .Y(N750) );
  AOI211X1TF U413 ( .A0(N546), .A1(N409), .B0(N752), .C0(N395), .Y(N761) );
  OAI21X1TF U414 ( .A0(N565), .A1(N233), .B0(N1151), .Y(N5000) );
  AOI22X1TF U415 ( .A0(N431), .A1(\GR[5][15] ), .B0(N432), .B1(\GR[7][15] ), 
        .Y(N1374) );
  OAI21X1TF U416 ( .A0(N569), .A1(N233), .B0(N1145), .Y(N4960) );
  AOI22X1TF U417 ( .A0(N341), .A1(\GR[5][11] ), .B0(N432), .B1(\GR[7][11] ), 
        .Y(N1358) );
  OAI21X1TF U418 ( .A0(N5750), .A1(N233), .B0(N1137), .Y(N490) );
  AOI22X1TF U419 ( .A0(N341), .A1(\GR[5][5] ), .B0(N1309), .B1(\GR[7][5] ), 
        .Y(N1334) );
  OAI21X1TF U420 ( .A0(N5760), .A1(N233), .B0(N1136), .Y(N489) );
  AOI22X1TF U421 ( .A0(N341), .A1(\GR[5][4] ), .B0(N1309), .B1(\GR[7][4] ), 
        .Y(N1330) );
  OAI21X1TF U422 ( .A0(N574), .A1(N233), .B0(N1139), .Y(N4910) );
  AOI22X1TF U423 ( .A0(N341), .A1(\GR[5][6] ), .B0(N1309), .B1(\GR[7][6] ), 
        .Y(N1338) );
  OAI21X1TF U424 ( .A0(N386), .A1(N227), .B0(N1098), .Y(N4700) );
  AOI22X1TF U425 ( .A0(N429), .A1(\GR[5][1] ), .B0(N430), .B1(\GR[7][1] ), .Y(
        N1246) );
  OAI21X1TF U426 ( .A0(N391), .A1(N227), .B0(N1113), .Y(N484) );
  AOI22X1TF U427 ( .A0(N342), .A1(\GR[5][15] ), .B0(N1237), .B1(\GR[7][15] ), 
        .Y(N1302) );
  OAI21X1TF U428 ( .A0(N397), .A1(N227), .B0(N1106), .Y(N478) );
  AOI22X1TF U429 ( .A0(N342), .A1(\GR[5][9] ), .B0(N1237), .B1(\GR[7][9] ), 
        .Y(N1278) );
  OAI21X1TF U430 ( .A0(N387), .A1(N227), .B0(N1102), .Y(N474) );
  AOI22X1TF U431 ( .A0(N429), .A1(\GR[5][5] ), .B0(N430), .B1(\GR[7][5] ), .Y(
        N1262) );
  OAI21X1TF U432 ( .A0(N379), .A1(N227), .B0(N1111), .Y(N483) );
  AOI22X1TF U433 ( .A0(N342), .A1(\GR[5][14] ), .B0(N1237), .B1(\GR[7][14] ), 
        .Y(N1298) );
  OAI21X1TF U434 ( .A0(N401), .A1(N227), .B0(N1110), .Y(N482) );
  AOI22X1TF U435 ( .A0(N342), .A1(\GR[5][13] ), .B0(N1237), .B1(\GR[7][13] ), 
        .Y(N1294) );
  OAI21X1TF U436 ( .A0(N402), .A1(N227), .B0(N1109), .Y(N481) );
  AOI22X1TF U437 ( .A0(N342), .A1(\GR[5][12] ), .B0(N1237), .B1(\GR[7][12] ), 
        .Y(N1290) );
  OAI21X1TF U438 ( .A0(N389), .A1(N227), .B0(N1100), .Y(N4720) );
  AOI22X1TF U439 ( .A0(N429), .A1(\GR[5][3] ), .B0(N430), .B1(\GR[7][3] ), .Y(
        N1254) );
  OAI21X1TF U440 ( .A0(N410), .A1(N228), .B0(N1108), .Y(N480) );
  AOI22X1TF U441 ( .A0(N342), .A1(\GR[5][11] ), .B0(N430), .B1(\GR[7][11] ), 
        .Y(N1286) );
  OAI21X1TF U442 ( .A0(N393), .A1(N228), .B0(N1101), .Y(N4730) );
  AOI22X1TF U443 ( .A0(N429), .A1(\GR[5][4] ), .B0(N430), .B1(\GR[7][4] ), .Y(
        N1258) );
  OAI21X1TF U444 ( .A0(N394), .A1(N228), .B0(N1099), .Y(N4710) );
  AOI22X1TF U445 ( .A0(N429), .A1(\GR[5][2] ), .B0(N430), .B1(\GR[7][2] ), .Y(
        N1250) );
  OAI21X1TF U446 ( .A0(N399), .A1(N228), .B0(N1104), .Y(N476) );
  AOI22X1TF U447 ( .A0(N429), .A1(\GR[5][7] ), .B0(N430), .B1(\GR[7][7] ), .Y(
        N1270) );
  OAI21X1TF U448 ( .A0(N400), .A1(N228), .B0(N1105), .Y(N477) );
  AOI22X1TF U449 ( .A0(N342), .A1(\GR[5][8] ), .B0(N1237), .B1(\GR[7][8] ), 
        .Y(N1274) );
  OAI21X1TF U450 ( .A0(N396), .A1(N228), .B0(N1103), .Y(N475) );
  AOI22X1TF U451 ( .A0(N429), .A1(\GR[5][6] ), .B0(N430), .B1(\GR[7][6] ), .Y(
        N1266) );
  OAI21X1TF U452 ( .A0(N411), .A1(N228), .B0(N1107), .Y(N479) );
  AOI22X1TF U453 ( .A0(N429), .A1(\GR[5][10] ), .B0(N430), .B1(\GR[7][10] ), 
        .Y(N1282) );
  OAI21X1TF U454 ( .A0(N392), .A1(N228), .B0(N1097), .Y(N4690) );
  AOI22X1TF U455 ( .A0(N429), .A1(\GR[5][0] ), .B0(N430), .B1(\GR[7][0] ), .Y(
        N1242) );
  AND3X2TF U456 ( .A(N94), .B(N92), .C(N93), .Y(N1237) );
  NOR3X1TF U457 ( .A(N93), .B(N382), .C(N376), .Y(N1236) );
  NOR3X4TF U458 ( .A(N92), .B(N93), .C(N376), .Y(N1234) );
  AND3X2TF U459 ( .A(N91), .B(N89), .C(N90), .Y(N1165) );
  NOR3X4TF U460 ( .A(N90), .B(N381), .C(N374), .Y(N1164) );
  OAI21X1TF U461 ( .A0(N1090), .A1(N1089), .B0(N1124), .Y(N1095) );
  OAI211X1TF U462 ( .A0(N1088), .A1(N1087), .B0(N1086), .C0(N1085), .Y(N1089)
         );
  OAI22X1TF U463 ( .A0(N390), .A1(N1094), .B0(N1120), .B1(N614), .Y(N1090) );
  OAI31X1TF U464 ( .A0(N755), .A1(CPU_WAIT), .A2(N754), .B0(N395), .Y(N756) );
  OAI21X1TF U465 ( .A0(N568), .A1(N233), .B0(N1146), .Y(N4970) );
  AOI22X1TF U466 ( .A0(N431), .A1(\GR[5][12] ), .B0(N432), .B1(\GR[7][12] ), 
        .Y(N1362) );
  OAI21X1TF U467 ( .A0(N570), .A1(N233), .B0(N1144), .Y(N4950) );
  AOI22X1TF U468 ( .A0(N431), .A1(\GR[5][10] ), .B0(N432), .B1(\GR[7][10] ), 
        .Y(N1354) );
  OAI21X1TF U469 ( .A0(N572), .A1(N234), .B0(N1142), .Y(N4930) );
  AOI22X1TF U470 ( .A0(N431), .A1(\GR[5][8] ), .B0(N432), .B1(\GR[7][8] ), .Y(
        N1346) );
  OAI21X1TF U471 ( .A0(N566), .A1(N234), .B0(N1149), .Y(N4990) );
  AOI22X1TF U472 ( .A0(N431), .A1(\GR[5][14] ), .B0(N432), .B1(\GR[7][14] ), 
        .Y(N1370) );
  OAI21X1TF U473 ( .A0(N571), .A1(N234), .B0(N1143), .Y(N4940) );
  AOI22X1TF U474 ( .A0(N431), .A1(\GR[5][9] ), .B0(N432), .B1(\GR[7][9] ), .Y(
        N1350) );
  OAI21X1TF U475 ( .A0(N567), .A1(N234), .B0(N1147), .Y(N4980) );
  AOI22X1TF U476 ( .A0(N431), .A1(\GR[5][13] ), .B0(N432), .B1(\GR[7][13] ), 
        .Y(N1366) );
  INVX2TF U477 ( .A(N1150), .Y(N1148) );
  OAI21X1TF U478 ( .A0(N573), .A1(N234), .B0(N1141), .Y(N4920) );
  AOI22X1TF U479 ( .A0(N431), .A1(\GR[5][7] ), .B0(N432), .B1(\GR[7][7] ), .Y(
        N1342) );
  OAI21X1TF U480 ( .A0(N371), .A1(N234), .B0(N1130), .Y(N485) );
  AOI22X1TF U481 ( .A0(N431), .A1(\GR[5][0] ), .B0(N1309), .B1(\GR[7][0] ), 
        .Y(N1314) );
  OAI21X1TF U482 ( .A0(N405), .A1(N234), .B0(N1132), .Y(N487) );
  AOI22X1TF U483 ( .A0(N341), .A1(\GR[5][2] ), .B0(N1309), .B1(\GR[7][2] ), 
        .Y(N1322) );
  AOI22X1TF U484 ( .A0(N341), .A1(\GR[5][1] ), .B0(N432), .B1(\GR[7][1] ), .Y(
        N1318) );
  OAI21X1TF U485 ( .A0(N1135), .A1(N2540), .B0(N1134), .Y(N488) );
  AOI22X1TF U486 ( .A0(N341), .A1(\GR[5][3] ), .B0(N1309), .B1(\GR[7][3] ), 
        .Y(N1326) );
  AND3X2TF U487 ( .A(N97), .B(N95), .C(N96), .Y(N1309) );
  NOR3X1TF U488 ( .A(N96), .B(N383), .C(N375), .Y(N1308) );
  NOR3X4TF U489 ( .A(N95), .B(N96), .C(N375), .Y(N1306) );
  INVX2TF U490 ( .A(N1133), .Y(N1135) );
  INVX2TF U491 ( .A(N1138), .Y(N1140) );
  NOR2X1TF U492 ( .A(N1128), .B(N1126), .Y(N1138) );
  AOI211X1TF U493 ( .A0(N22), .A1(N1123), .B0(N1122), .C0(N1121), .Y(N1126) );
  INVX2TF U494 ( .A(N1040), .Y(N600) );
  AOI21X1TF U495 ( .A0(N975), .A1(N1087), .B0(N1088), .Y(N1118) );
  OAI22X1TF U496 ( .A0(N746), .A1(N423), .B0(N745), .B1(N744), .Y(N747) );
  OAI21X1TF U497 ( .A0(N743), .A1(I_ADDR[8]), .B0(N742), .Y(N744) );
  OAI22X1TF U498 ( .A0(N746), .A1(N420), .B0(N745), .B1(N737), .Y(N738) );
  OAI22X1TF U499 ( .A0(N746), .A1(N421), .B0(N745), .B1(N725), .Y(N726) );
  OAI22X1TF U500 ( .A0(N746), .A1(N422), .B0(N745), .B1(N731), .Y(N732) );
  NOR2X1TF U501 ( .A(N746), .B(N415), .Y(N740) );
  AOI211X1TF U502 ( .A0(N739), .A1(N415), .B0(N743), .C0(N745), .Y(N741) );
  NOR2X1TF U503 ( .A(N746), .B(N417), .Y(N656) );
  AOI211X1TF U504 ( .A0(N742), .A1(N417), .B0(N882), .C0(N745), .Y(N657) );
  NOR2X1TF U505 ( .A(N742), .B(N417), .Y(N882) );
  NOR2X1TF U506 ( .A(N739), .B(N415), .Y(N743) );
  NOR2X1TF U507 ( .A(N746), .B(N414), .Y(N734) );
  AOI211X1TF U508 ( .A0(N733), .A1(N414), .B0(N736), .C0(N745), .Y(N735) );
  NOR2X1TF U509 ( .A(N733), .B(N414), .Y(N736) );
  AOI22X1TF U510 ( .A0(I_ADDR[1]), .A1(N746), .B0(N745), .B1(N419), .Y(N655)
         );
  NOR2X1TF U511 ( .A(N746), .B(N413), .Y(N728) );
  AOI211X1TF U512 ( .A0(N727), .A1(N413), .B0(N730), .C0(N745), .Y(N729) );
  NAND3X2TF U513 ( .A(N670), .B(N654), .C(N746), .Y(N745) );
  OAI211X4TF U514 ( .A0(N659), .A1(N653), .B0(N751), .C0(N345), .Y(N746) );
  OR2X2TF U515 ( .A(INSTR_OVER), .B(N690), .Y(N751) );
  NOR2X1TF U516 ( .A(N727), .B(N413), .Y(N730) );
  AOI32X1TF U517 ( .A0(N652), .A1(N1122), .A2(N651), .B0(N650), .B1(N1122), 
        .Y(N654) );
  AOI21X1TF U518 ( .A0(N606), .A1(ZF), .B0(N649), .Y(N652) );
  AOI22X1TF U519 ( .A0(N335), .A1(N1157), .B0(N560), .B1(N1156), .Y(N517) );
  AOI22X1TF U520 ( .A0(N2200), .A1(N1155), .B0(N2550), .B1(N1153), .Y(N5010)
         );
  AOI22X1TF U521 ( .A0(N2200), .A1(N1157), .B0(N2540), .B1(N1153), .Y(N5050)
         );
  INVX2TF U522 ( .A(I_DATAIN[3]), .Y(N1157) );
  AOI22X1TF U523 ( .A0(N335), .A1(N1155), .B0(N384), .B1(N1156), .Y(N513) );
  INVX2TF U524 ( .A(I_DATAIN[7]), .Y(N1155) );
  INVX2TF U525 ( .A(N606), .Y(N975) );
  NOR2X1TF U526 ( .A(N599), .B(N661), .Y(N959) );
  INVX2TF U527 ( .A(N1124), .Y(N1128) );
  OAI211X1TF U528 ( .A0(N546), .A1(N659), .B0(N668), .C0(N424), .Y(N748) );
  INVX2TF U529 ( .A(N749), .Y(N659) );
  NOR3X1TF U530 ( .A(N409), .B(STATE[3]), .C(STATE[1]), .Y(N749) );
  AOI22X2TF U531 ( .A0(D_ADDR[9]), .A1(N692), .B0(N694), .B1(D_DATAIN[0]), .Y(
        N709) );
  AOI22X2TF U532 ( .A0(D_ADDR[2]), .A1(N670), .B0(N669), .B1(D_DATAIN[1]), .Y(
        N682) );
  AOI22X2TF U533 ( .A0(D_ADDR[1]), .A1(N670), .B0(N669), .B1(D_DATAIN[0]), .Y(
        N681) );
  AOI22X2TF U534 ( .A0(D_ADDR[5]), .A1(N670), .B0(N669), .B1(D_DATAIN[4]), .Y(
        N685) );
  AOI22X2TF U535 ( .A0(D_ADDR[8]), .A1(N670), .B0(N669), .B1(D_DATAIN[7]), .Y(
        N688) );
  AOI22X2TF U536 ( .A0(D_ADDR[6]), .A1(N670), .B0(N669), .B1(D_DATAIN[5]), .Y(
        N686) );
  AOI22X2TF U537 ( .A0(D_ADDR[3]), .A1(N670), .B0(N669), .B1(D_DATAIN[2]), .Y(
        N683) );
  AOI22X2TF U538 ( .A0(D_ADDR[7]), .A1(N670), .B0(N669), .B1(D_DATAIN[6]), .Y(
        N687) );
  AOI22X2TF U539 ( .A0(D_ADDR[4]), .A1(N670), .B0(N669), .B1(D_DATAIN[3]), .Y(
        N684) );
  AOI32X4TF U540 ( .A0(N667), .A1(N691), .A2(N612), .B0(N666), .B1(N691), .Y(
        N693) );
  OAI211X1TF U541 ( .A0(N1116), .A1(N665), .B0(N664), .C0(N663), .Y(N666) );
  OAI211X1TF U542 ( .A0(N597), .A1(N199), .B0(N1060), .C0(N1059), .Y(N388) );
  AOI22X1TF U543 ( .A0(IO_DATAINB[5]), .A1(N334), .B0(N1081), .B1(N1058), .Y(
        N1059) );
  AOI22X1TF U544 ( .A0(IO_DATAINA[5]), .A1(N2150), .B0(D_ADDR[6]), .B1(N1079), 
        .Y(N1060) );
  OAI211X1TF U545 ( .A0(N1063), .A1(N331), .B0(N1055), .C0(N1054), .Y(N358) );
  AOI22X1TF U546 ( .A0(IO_DATAINB[12]), .A1(N593), .B0(N1075), .B1(N1053), .Y(
        N1054) );
  INVX2TF U547 ( .A(N605), .Y(N1053) );
  OAI211X1TF U548 ( .A0(N1063), .A1(N199), .B0(N1062), .C0(N1061), .Y(N398) );
  AOI22X1TF U549 ( .A0(IO_DATAINB[11]), .A1(N334), .B0(N1081), .B1(N1064), .Y(
        N1061) );
  NOR4X1TF U550 ( .A(N1039), .B(N1038), .C(N1037), .D(N1036), .Y(N1063) );
  OAI22X1TF U551 ( .A0(N511), .A1(N410), .B0(N1035), .B1(N1034), .Y(N512) );
  AOI21X1TF U552 ( .A0(N433), .A1(N569), .B0(N201), .Y(N511) );
  OAI22X1TF U553 ( .A0(N1030), .A1(N1029), .B0(N1028), .B1(N1027), .Y(N1037)
         );
  INVX2TF U554 ( .A(N1026), .Y(N1030) );
  AOI21X1TF U555 ( .A0(N615), .A1(N1022), .B0(N569), .Y(N1039) );
  AOI22X1TF U556 ( .A0(REG_A[11]), .A1(N610), .B0(N434), .B1(N410), .Y(N1022)
         );
  OAI211X1TF U557 ( .A0(N598), .A1(N331), .B0(N1049), .C0(N1048), .Y(N338) );
  AOI22X1TF U558 ( .A0(IO_DATAINB[8]), .A1(N334), .B0(N1075), .B1(N1050), .Y(
        N1048) );
  AOI22X1TF U559 ( .A0(IO_DATAINA[8]), .A1(N2150), .B0(D_ADDR[9]), .B1(N1079), 
        .Y(N1049) );
  OAI211X1TF U560 ( .A0(N598), .A1(N199), .B0(N1083), .C0(N1082), .Y(N4680) );
  AOI22X1TF U561 ( .A0(IO_DATAINB[7]), .A1(N334), .B0(N1081), .B1(N1080), .Y(
        N1082) );
  AOI22X1TF U562 ( .A0(IO_DATAINA[7]), .A1(N2150), .B0(D_ADDR[8]), .B1(N1079), 
        .Y(N1083) );
  AOI211X1TF U563 ( .A0(N498), .A1(N280), .B0(N555), .C0(N554), .Y(N598) );
  AOI211X1TF U564 ( .A0(N604), .A1(N1026), .B0(N981), .C0(N980), .Y(N982) );
  OAI21X1TF U565 ( .A0(N979), .A1(N1027), .B0(N978), .Y(N980) );
  OAI22X1TF U566 ( .A0(N1025), .A1(N1028), .B0(N976), .B1(N399), .Y(N981) );
  AOI21X1TF U567 ( .A0(N434), .A1(N573), .B0(N201), .Y(N976) );
  AOI21X1TF U568 ( .A0(N615), .A1(N553), .B0(N573), .Y(N555) );
  AOI22X1TF U569 ( .A0(N610), .A1(REG_A[7]), .B0(N433), .B1(N399), .Y(N553) );
  OAI211X1TF U570 ( .A0(N597), .A1(N331), .B0(N1077), .C0(N1076), .Y(N4580) );
  AOI22X1TF U571 ( .A0(IO_DATAINB[6]), .A1(N334), .B0(N1075), .B1(N1080), .Y(
        N1076) );
  AOI22X1TF U572 ( .A0(IO_DATAINA[6]), .A1(N2150), .B0(D_ADDR[7]), .B1(N1079), 
        .Y(N1077) );
  AND3X2TF U573 ( .A(N582), .B(N782), .C(N581), .Y(N597) );
  AOI211X1TF U574 ( .A0(N1018), .A1(N1010), .B0(N781), .C0(N780), .Y(N782) );
  OAI22X1TF U575 ( .A0(N779), .A1(N995), .B0(N985), .B1(N979), .Y(N780) );
  AOI21X1TF U576 ( .A0(N434), .A1(N5750), .B0(N201), .Y(N778) );
  AOI22X1TF U577 ( .A0(N344), .A1(REG_A[5]), .B0(N433), .B1(N387), .Y(N579) );
  AOI22X1TF U578 ( .A0(N2160), .A1(IO_DATAINA[1]), .B0(N334), .B1(
        IO_DATAINB[1]), .Y(N1046) );
  AOI22X1TF U579 ( .A0(IO_STATUS[1]), .A1(N595), .B0(D_ADDR[2]), .B1(N1079), 
        .Y(N1047) );
  OAI211X1TF U580 ( .A0(N1067), .A1(N331), .B0(N1066), .C0(N1065), .Y(N408) );
  AOI22X1TF U581 ( .A0(IO_DATAINB[10]), .A1(N334), .B0(N1075), .B1(N1064), .Y(
        N1065) );
  OAI211X1TF U582 ( .A0(N1067), .A1(N199), .B0(N1052), .C0(N1051), .Y(N348) );
  AOI22X1TF U583 ( .A0(IO_DATAINB[9]), .A1(N334), .B0(N1081), .B1(N1050), .Y(
        N1051) );
  INVX2TF U584 ( .A(N583), .Y(N1050) );
  AOI211X1TF U585 ( .A0(N499), .A1(N279), .B0(N538), .C0(N537), .Y(N583) );
  AOI211X1TF U586 ( .A0(N604), .A1(N963), .B0(N962), .C0(N961), .Y(N964) );
  OAI21X1TF U587 ( .A0(N1029), .A1(N830), .B0(N829), .Y(N961) );
  OAI22X1TF U588 ( .A0(N827), .A1(N1028), .B0(N826), .B1(N400), .Y(N962) );
  AOI21X1TF U589 ( .A0(N434), .A1(N572), .B0(N201), .Y(N826) );
  AOI21X1TF U590 ( .A0(N615), .A1(N536), .B0(N572), .Y(N538) );
  AOI22X1TF U591 ( .A0(N610), .A1(REG_A[8]), .B0(N433), .B1(N400), .Y(N536) );
  AOI211X1TF U592 ( .A0(N604), .A1(N1021), .B0(N1020), .C0(N1019), .Y(N1067)
         );
  AOI211X1TF U593 ( .A0(N466), .A1(N425), .B0(N4670), .C0(N385), .Y(N510) );
  AOI21X1TF U594 ( .A0(N615), .A1(N4660), .B0(N571), .Y(N4670) );
  AOI22X1TF U595 ( .A0(N610), .A1(REG_A[9]), .B0(N433), .B1(N397), .Y(N4660)
         );
  OAI31X1TF U596 ( .A0(N407), .A1(N1014), .A2(N1013), .B0(N1012), .Y(N1020) );
  OAI211X1TF U597 ( .A0(N1070), .A1(N1078), .B0(N1069), .C0(N1068), .Y(N1071)
         );
  AOI22X1TF U598 ( .A0(N2150), .A1(IO_DATAINA[2]), .B0(N595), .B1(IO_STATUS[2]), .Y(N1068) );
  AOI22X1TF U599 ( .A0(IO_DATAINB[2]), .A1(N593), .B0(D_ADDR[3]), .B1(N424), 
        .Y(N1069) );
  AOI211X1TF U600 ( .A0(REG_B[1]), .A1(N1002), .B0(N1001), .C0(N1000), .Y(
        N1070) );
  OAI211X1TF U601 ( .A0(N998), .A1(N999), .B0(N997), .C0(N4650), .Y(N1000) );
  AOI22X1TF U602 ( .A0(N279), .A1(N492), .B0(N458), .B1(N425), .Y(N4650) );
  OAI211X1TF U603 ( .A0(N393), .A1(N332), .B0(N992), .C0(N991), .Y(N996) );
  INVX2TF U604 ( .A(N985), .Y(N1017) );
  NOR2X1TF U605 ( .A(N804), .B(N387), .Y(N777) );
  OAI32X1TF U606 ( .A0(N386), .A1(REG_B[1]), .A2(N373), .B0(N984), .B1(N386), 
        .Y(N1001) );
  OAI211X1TF U607 ( .A0(N596), .A1(N331), .B0(N1057), .C0(N1056), .Y(N378) );
  AOI22X1TF U608 ( .A0(IO_DATAINB[4]), .A1(N334), .B0(N1075), .B1(N1058), .Y(
        N1056) );
  OR4X2TF U609 ( .A(N535), .B(N825), .C(N824), .D(N534), .Y(N1058) );
  OAI21X1TF U610 ( .A0(N1034), .A1(N830), .B0(N823), .Y(N824) );
  INVX2TF U611 ( .A(N965), .Y(N827) );
  INVX2TF U612 ( .A(N818), .Y(N830) );
  INVX2TF U613 ( .A(N604), .Y(N1034) );
  AOI21X1TF U614 ( .A0(N435), .A1(N5760), .B0(N201), .Y(N817) );
  AOI21X1TF U615 ( .A0(N615), .A1(N532), .B0(N5760), .Y(N535) );
  AOI22X1TF U616 ( .A0(N344), .A1(REG_A[4]), .B0(N433), .B1(N393), .Y(N532) );
  INVX2TF U617 ( .A(N198), .Y(N1075) );
  AOI22X1TF U618 ( .A0(IO_DATAINA[4]), .A1(N2160), .B0(D_ADDR[5]), .B1(N1079), 
        .Y(N1057) );
  OAI211X1TF U619 ( .A0(N596), .A1(N199), .B0(N1074), .C0(N1073), .Y(N428) );
  AOI22X1TF U620 ( .A0(IO_DATAINB[3]), .A1(N334), .B0(N1081), .B1(N1072), .Y(
        N1073) );
  AOI211X1TF U621 ( .A0(N493), .A1(N280), .B0(N795), .C0(N529), .Y(N531) );
  INVX2TF U622 ( .A(N785), .Y(N796) );
  OAI211X1TF U623 ( .A0(N393), .A1(N969), .B0(N784), .C0(N783), .Y(N785) );
  OAI22X1TF U624 ( .A0(N1003), .A1(N608), .B0(N1005), .B1(N791), .Y(N795) );
  OAI22X1TF U625 ( .A0(N793), .A1(N394), .B0(N792), .B1(N197), .Y(N794) );
  AOI221X1TF U626 ( .A0(N434), .A1(N394), .B0(N610), .B1(REG_A[2]), .C0(N1015), 
        .Y(N792) );
  INVX2TF U627 ( .A(N1078), .Y(N1081) );
  AOI22X1TF U628 ( .A0(IO_DATAINA[3]), .A1(N2150), .B0(D_ADDR[4]), .B1(N1079), 
        .Y(N1074) );
  AND3X2TF U629 ( .A(N811), .B(N812), .C(N558), .Y(N596) );
  AOI21X1TF U630 ( .A0(N1026), .A1(N2140), .B0(N557), .Y(N558) );
  AOI22X1TF U631 ( .A0(N799), .A1(N616), .B0(N460), .B1(N425), .Y(N556) );
  OAI211X1TF U632 ( .A0(N332), .A1(N396), .B0(N798), .C0(N797), .Y(N799) );
  AOI211X1TF U633 ( .A0(REG_A[14]), .A1(N807), .B0(N806), .C0(N805), .Y(N1025)
         );
  OAI22X1TF U634 ( .A0(N401), .A1(N969), .B0(N410), .B1(N804), .Y(N806) );
  INVX2TF U635 ( .A(N1028), .Y(N1018) );
  AOI221X1TF U636 ( .A0(N389), .A1(N434), .B0(REG_A[3]), .B1(N344), .C0(N808), 
        .Y(N809) );
  OAI31X1TF U637 ( .A0(N998), .A1(N197), .A2(N1027), .B0(N615), .Y(N808) );
  OAI21X1TF U638 ( .A0(REG_B[3]), .A1(N373), .B0(N984), .Y(N810) );
  OAI211X1TF U639 ( .A0(N637), .A1(N1014), .B0(N4630), .C0(N4620), .Y(N4640)
         );
  AOI211X1TF U640 ( .A0(N634), .A1(N2140), .B0(N4610), .C0(N4600), .Y(N4620)
         );
  OAI22X1TF U641 ( .A0(N768), .A1(N1004), .B0(N566), .B1(N638), .Y(N4600) );
  AOI221X1TF U642 ( .A0(N434), .A1(N379), .B0(N610), .B1(REG_A[14]), .C0(N1015), .Y(N638) );
  NOR2X1TF U643 ( .A(N4590), .B(N379), .Y(N4610) );
  AOI21X1TF U644 ( .A0(N433), .A1(N566), .B0(N643), .Y(N4590) );
  OAI211X1TF U645 ( .A0(N332), .A1(N410), .B0(N633), .C0(N632), .Y(N634) );
  AOI21X1TF U646 ( .A0(IO_DATAINA[0]), .A1(N2160), .B0(N589), .Y(N590) );
  OAI211X1TF U647 ( .A0(N601), .A1(N198), .B0(N588), .C0(N587), .Y(N589) );
  AOI22X1TF U648 ( .A0(N593), .A1(IO_DATAINB[0]), .B0(D_ADDR[1]), .B1(N424), 
        .Y(N588) );
  NOR2X1TF U649 ( .A(N663), .B(N452), .Y(N453) );
  AND2X2TF U650 ( .A(N560), .B(N384), .Y(N452) );
  OAI211X1TF U651 ( .A0(N998), .A1(N974), .B0(N973), .C0(N564), .Y(N577) );
  AOI21X1TF U652 ( .A0(N279), .A1(N491), .B0(N563), .Y(N564) );
  OAI21X1TF U653 ( .A0(REG_B[0]), .A1(N373), .B0(N561), .Y(N562) );
  OAI31X1TF U654 ( .A0(N972), .A1(N971), .A2(N970), .B0(N616), .Y(N973) );
  NOR2X1TF U655 ( .A(N969), .B(N394), .Y(N970) );
  NOR2X1TF U656 ( .A(N968), .B(N386), .Y(N972) );
  NOR2X1TF U657 ( .A(N993), .B(N410), .Y(N816) );
  INVX2TF U658 ( .A(N790), .Y(N998) );
  OAI211X1TF U659 ( .A0(REG_A[0]), .A1(N436), .B0(N615), .C0(N559), .Y(N578)
         );
  INVX2TF U660 ( .A(N612), .Y(N1088) );
  INVX2TF U661 ( .A(N1043), .Y(N1064) );
  AND2X2TF U662 ( .A(N528), .B(N527), .Y(N1043) );
  AOI21X1TF U663 ( .A0(N467), .A1(N425), .B0(N526), .Y(N527) );
  NOR2X1TF U664 ( .A(N1008), .B(N523), .Y(N524) );
  AOI22X1TF U665 ( .A0(N1006), .A1(N2130), .B0(REG_A[10]), .B1(N1007), .Y(N522) );
  NOR2X1TF U666 ( .A(N993), .B(N389), .Y(N971) );
  OAI22X1TF U667 ( .A0(N1005), .A1(N1004), .B0(N1003), .B1(N1029), .Y(N1008)
         );
  INVX2TF U668 ( .A(N787), .Y(N1003) );
  OAI21X1TF U669 ( .A0(N969), .A1(N392), .B0(N636), .Y(N787) );
  AOI22X1TF U670 ( .A0(N641), .A1(REG_A[1]), .B0(N2210), .B1(REG_A[2]), .Y(
        N636) );
  AOI22X1TF U671 ( .A0(REG_B[2]), .A1(N789), .B0(N788), .B1(N197), .Y(N1005)
         );
  OAI211X1TF U672 ( .A0(N411), .A1(N804), .B0(N763), .C0(N762), .Y(N788) );
  AOI22X1TF U673 ( .A0(REG_A[13]), .A1(N807), .B0(REG_A[12]), .B1(N426), .Y(
        N762) );
  AOI221X1TF U674 ( .A0(REG_B[0]), .A1(N391), .B0(N371), .B1(N379), .C0(
        REG_B[1]), .Y(N789) );
  AND2X2TF U675 ( .A(N450), .B(N449), .Y(N605) );
  AOI21X1TF U676 ( .A0(N469), .A1(N425), .B0(N447), .Y(N449) );
  OAI211X1TF U677 ( .A0(N993), .A1(N397), .B0(N763), .C0(N814), .Y(N618) );
  OAI211X1TF U678 ( .A0(N391), .A1(N993), .B0(N617), .C0(N632), .Y(N965) );
  AOI22X1TF U679 ( .A0(REG_A[12]), .A1(N2220), .B0(N426), .B1(REG_A[14]), .Y(
        N617) );
  AOI221X1TF U680 ( .A0(N434), .A1(N402), .B0(N610), .B1(REG_A[12]), .C0(N1015), .Y(N622) );
  OAI211X1TF U681 ( .A0(N386), .A1(N993), .B0(N620), .C0(N784), .Y(N963) );
  AOI22X1TF U682 ( .A0(N426), .A1(REG_A[2]), .B0(N2210), .B1(REG_A[4]), .Y(
        N620) );
  NOR2X1TF U683 ( .A(N804), .B(N392), .Y(N818) );
  NOR3X1TF U684 ( .A(N630), .B(N631), .C(N455), .Y(N456) );
  AOI211X1TF U685 ( .A0(N343), .A1(REG_A[11]), .B0(N803), .C0(N805), .Y(N454)
         );
  NOR2X1TF U686 ( .A(N402), .B(N968), .Y(N805) );
  NOR2X1TF U687 ( .A(N993), .B(N411), .Y(N803) );
  OAI22X1TF U688 ( .A0(N779), .A1(N627), .B0(N985), .B1(N1024), .Y(N631) );
  AOI21X1TF U689 ( .A0(REG_A[13]), .A1(N2210), .B0(N626), .Y(N985) );
  OAI22X1TF U690 ( .A0(N969), .A1(N391), .B0(N968), .B1(N379), .Y(N626) );
  OAI211X1TF U691 ( .A0(N394), .A1(N993), .B0(N625), .C0(N798), .Y(N1021) );
  AOI22X1TF U692 ( .A0(N343), .A1(REG_A[3]), .B0(N2220), .B1(REG_A[5]), .Y(
        N625) );
  OAI22X1TF U693 ( .A0(N567), .A1(N629), .B0(N628), .B1(N401), .Y(N630) );
  AOI21X1TF U694 ( .A0(N435), .A1(N567), .B0(N643), .Y(N628) );
  INVX2TF U695 ( .A(N436), .Y(N435) );
  AOI221X1TF U696 ( .A0(N434), .A1(N401), .B0(N610), .B1(REG_A[13]), .C0(N1015), .Y(N629) );
  INVX2TF U697 ( .A(N436), .Y(N434) );
  OAI211X1TF U698 ( .A0(N565), .A1(N551), .B0(N550), .C0(N549), .Y(N552) );
  AOI211X1TF U699 ( .A0(N604), .A1(N1023), .B0(N548), .C0(N547), .Y(N549) );
  OAI21X1TF U700 ( .A0(N544), .A1(N391), .B0(N543), .Y(N547) );
  OAI22X1TF U701 ( .A0(N969), .A1(N401), .B0(N968), .B1(N379), .Y(N542) );
  INVX2TF U702 ( .A(N426), .Y(N969) );
  NOR2X1TF U703 ( .A(N993), .B(N402), .Y(N771) );
  AOI21X1TF U704 ( .A0(N565), .A1(N433), .B0(N541), .Y(N544) );
  NOR2X2TF U705 ( .A(N1044), .B(N1127), .Y(N790) );
  INVX2TF U706 ( .A(N436), .Y(N433) );
  NOR2X1TF U707 ( .A(N540), .B(N1014), .Y(N548) );
  INVX2TF U708 ( .A(N609), .Y(N1014) );
  NOR2X2TF U709 ( .A(REG_B[2]), .B(N407), .Y(N986) );
  NOR2X1TF U710 ( .A(N407), .B(N197), .Y(N987) );
  OAI211X1TF U711 ( .A0(N392), .A1(N993), .B0(N642), .C0(N991), .Y(N1026) );
  AOI22X1TF U712 ( .A0(N343), .A1(REG_A[1]), .B0(N2220), .B1(REG_A[3]), .Y(
        N642) );
  NOR2X1TF U713 ( .A(N406), .B(REG_B[0]), .Y(N990) );
  INVX2TF U714 ( .A(N968), .Y(N641) );
  AND2X2TF U715 ( .A(N609), .B(N988), .Y(N604) );
  AND2X2TF U716 ( .A(N1086), .B(N439), .Y(N440) );
  NOR2X1TF U717 ( .A(CODE_TYPE[1]), .B(N560), .Y(N619) );
  AOI211X1TF U718 ( .A0(N344), .A1(REG_A[15]), .B0(N1015), .C0(N539), .Y(N551)
         );
  NOR2X1TF U719 ( .A(N373), .B(REG_A[15]), .Y(N539) );
  NAND2X2TF U720 ( .A(N613), .B(N1123), .Y(N373) );
  AOI211X1TF U721 ( .A0(N612), .A1(N1123), .B0(N611), .C0(N200), .Y(N647) );
  INVX2TF U722 ( .A(N1091), .Y(N1116) );
  OR2X2TF U723 ( .A(N1125), .B(N665), .Y(N983) );
  INVX2TF U724 ( .A(N613), .Y(N665) );
  OAI21X1TF U725 ( .A0(N1042), .A1(N1115), .B0(N613), .Y(N437) );
  NOR2BX2TF U726 ( .AN(CODE_TYPE[3]), .B(N2100), .Y(N613) );
  AOI22X1TF U727 ( .A0(N1306), .A1(N1389), .B0(N291), .B1(\GR[6][15] ), .Y(
        N1373) );
  AOI22X1TF U728 ( .A0(N313), .A1(N1375), .B0(N273), .B1(N1386), .Y(N1372) );
  AOI22X1TF U729 ( .A0(N315), .A1(\GR[0][15] ), .B0(N277), .B1(N1383), .Y(
        N1371) );
  AOI22X1TF U730 ( .A0(N350), .A1(N1393), .B0(N290), .B1(\GR[6][11] ), .Y(
        N1357) );
  AOI22X1TF U731 ( .A0(N313), .A1(N1379), .B0(N273), .B1(N35), .Y(N1356) );
  AOI22X1TF U732 ( .A0(N315), .A1(\GR[0][11] ), .B0(N277), .B1(IO_DATAOUTA[11]), .Y(N1355) );
  AOI22X1TF U733 ( .A0(N224), .A1(N257), .B0(N1138), .B1(N93), .Y(N1137) );
  AOI22X1TF U734 ( .A0(N350), .A1(IO_OFFSET[5]), .B0(N291), .B1(\GR[6][5] ), 
        .Y(N1333) );
  AOI22X1TF U735 ( .A0(N315), .A1(\GR[0][5] ), .B0(N277), .B1(IO_DATAOUTA[5]), 
        .Y(N1331) );
  AOI22X1TF U736 ( .A0(N224), .A1(N258), .B0(N1138), .B1(N92), .Y(N1136) );
  AOI22X1TF U737 ( .A0(N350), .A1(IO_OFFSET[4]), .B0(N291), .B1(\GR[6][4] ), 
        .Y(N1329) );
  AOI22X1TF U738 ( .A0(N313), .A1(\IO_CONTROL[4] ), .B0(N273), .B1(N30), .Y(
        N1328) );
  AOI22X1TF U739 ( .A0(N315), .A1(\GR[0][4] ), .B0(N277), .B1(N26), .Y(N1327)
         );
  AOI22X1TF U740 ( .A0(N224), .A1(N256), .B0(N1138), .B1(N94), .Y(N1139) );
  AOI22X1TF U741 ( .A0(N350), .A1(IO_OFFSET[6]), .B0(N291), .B1(\GR[6][6] ), 
        .Y(N1337) );
  AOI22X1TF U742 ( .A0(N315), .A1(\GR[0][6] ), .B0(N277), .B1(N27), .Y(N1335)
         );
  AOI22X1TF U743 ( .A0(N310), .A1(\IO_CONTROL[1] ), .B0(N268), .B1(
        IO_DATAOUTB[1]), .Y(N1244) );
  AOI22X1TF U744 ( .A0(N316), .A1(\GR[0][1] ), .B0(N274), .B1(N24), .Y(N1243)
         );
  AOI22X1TF U745 ( .A0(N1164), .A1(\GR[5][1] ), .B0(N427), .B1(\GR[7][1] ), 
        .Y(N1174) );
  AOI22X1TF U746 ( .A0(N292), .A1(\IO_CONTROL[1] ), .B0(N270), .B1(
        IO_DATAOUTB[1]), .Y(N1172) );
  AOI22X1TF U747 ( .A0(N310), .A1(N1375), .B0(N268), .B1(N1386), .Y(N1300) );
  AOI22X1TF U748 ( .A0(N316), .A1(\GR[0][15] ), .B0(N274), .B1(N1383), .Y(
        N1299) );
  AOI22X1TF U749 ( .A0(N1164), .A1(\GR[5][15] ), .B0(N1165), .B1(\GR[7][15] ), 
        .Y(N1230) );
  AOI22X1TF U750 ( .A0(N232), .A1(N1389), .B0(N282), .B1(\GR[6][15] ), .Y(
        N1229) );
  AOI22X1TF U751 ( .A0(N309), .A1(N1375), .B0(N271), .B1(N1386), .Y(N1228) );
  AOI22X1TF U752 ( .A0(N230), .A1(\GR[0][15] ), .B0(N284), .B1(N1383), .Y(
        N1227) );
  AOI22X1TF U753 ( .A0(N310), .A1(N1381), .B0(N268), .B1(IO_DATAOUTB[9]), .Y(
        N1276) );
  AOI22X1TF U754 ( .A0(N316), .A1(\GR[0][9] ), .B0(N274), .B1(N32), .Y(N1275)
         );
  AOI22X1TF U755 ( .A0(N1164), .A1(\GR[5][9] ), .B0(N1165), .B1(\GR[7][9] ), 
        .Y(N1206) );
  AOI22X1TF U756 ( .A0(N232), .A1(IO_OFFSET[9]), .B0(N282), .B1(\GR[6][9] ), 
        .Y(N1205) );
  AOI22X1TF U757 ( .A0(N309), .A1(N1381), .B0(N271), .B1(IO_DATAOUTB[9]), .Y(
        N1204) );
  AOI22X1TF U758 ( .A0(N230), .A1(\GR[0][9] ), .B0(N284), .B1(N32), .Y(N1203)
         );
  AOI22X1TF U759 ( .A0(N316), .A1(\GR[0][5] ), .B0(N274), .B1(IO_DATAOUTA[5]), 
        .Y(N1259) );
  AOI22X1TF U760 ( .A0(N1164), .A1(\GR[5][5] ), .B0(N427), .B1(\GR[7][5] ), 
        .Y(N1190) );
  AOI22X1TF U761 ( .A0(N311), .A1(N1376), .B0(N268), .B1(N1387), .Y(N1296) );
  AOI22X1TF U762 ( .A0(N317), .A1(\GR[0][14] ), .B0(N274), .B1(N1384), .Y(
        N1295) );
  AOI22X1TF U763 ( .A0(N1164), .A1(\GR[5][14] ), .B0(N1165), .B1(\GR[7][14] ), 
        .Y(N1226) );
  AOI22X1TF U764 ( .A0(N232), .A1(N1390), .B0(N282), .B1(\GR[6][14] ), .Y(
        N1225) );
  AOI22X1TF U765 ( .A0(N309), .A1(N1376), .B0(N271), .B1(N1387), .Y(N1224) );
  AOI22X1TF U766 ( .A0(N230), .A1(\GR[0][14] ), .B0(N284), .B1(N1384), .Y(
        N1223) );
  AOI22X1TF U767 ( .A0(N1234), .A1(N1391), .B0(N286), .B1(\GR[6][13] ), .Y(
        N1293) );
  AOI22X1TF U768 ( .A0(N311), .A1(N1377), .B0(N269), .B1(N1388), .Y(N1292) );
  AOI22X1TF U769 ( .A0(N317), .A1(\GR[0][13] ), .B0(N275), .B1(N1385), .Y(
        N1291) );
  AOI22X1TF U770 ( .A0(N1164), .A1(\GR[5][13] ), .B0(N1165), .B1(\GR[7][13] ), 
        .Y(N1222) );
  AOI22X1TF U771 ( .A0(N232), .A1(N1391), .B0(N282), .B1(\GR[6][13] ), .Y(
        N1221) );
  AOI22X1TF U772 ( .A0(N309), .A1(N1377), .B0(N271), .B1(N1388), .Y(N1220) );
  AOI22X1TF U773 ( .A0(N230), .A1(\GR[0][13] ), .B0(N284), .B1(N1385), .Y(
        N1219) );
  AOI22X1TF U774 ( .A0(N1234), .A1(N1392), .B0(N286), .B1(\GR[6][12] ), .Y(
        N1289) );
  AOI22X1TF U775 ( .A0(N311), .A1(N1378), .B0(N269), .B1(IO_DATAOUTB[12]), .Y(
        N1288) );
  AOI22X1TF U776 ( .A0(N317), .A1(\GR[0][12] ), .B0(N275), .B1(N34), .Y(N1287)
         );
  AOI22X1TF U777 ( .A0(N1164), .A1(\GR[5][12] ), .B0(N1165), .B1(\GR[7][12] ), 
        .Y(N1218) );
  AOI22X1TF U778 ( .A0(N292), .A1(N1378), .B0(N270), .B1(IO_DATAOUTB[12]), .Y(
        N1216) );
  AOI22X1TF U779 ( .A0(N351), .A1(IO_OFFSET[3]), .B0(N286), .B1(\GR[6][3] ), 
        .Y(N1253) );
  AOI22X1TF U780 ( .A0(N311), .A1(\IO_CONTROL[3] ), .B0(N269), .B1(N29), .Y(
        N1252) );
  AOI22X1TF U781 ( .A0(N317), .A1(\GR[0][3] ), .B0(N275), .B1(IO_DATAOUTA[3]), 
        .Y(N1251) );
  AOI22X1TF U782 ( .A0(N1164), .A1(\GR[5][3] ), .B0(N427), .B1(\GR[7][3] ), 
        .Y(N1182) );
  AOI22X1TF U783 ( .A0(N232), .A1(IO_OFFSET[3]), .B0(N282), .B1(\GR[6][3] ), 
        .Y(N1181) );
  AOI22X1TF U784 ( .A0(N309), .A1(\IO_CONTROL[3] ), .B0(N271), .B1(N29), .Y(
        N1180) );
  AOI22X1TF U785 ( .A0(N230), .A1(\GR[0][3] ), .B0(N284), .B1(IO_DATAOUTA[3]), 
        .Y(N1179) );
  AOI22X1TF U786 ( .A0(N351), .A1(N1393), .B0(N286), .B1(\GR[6][11] ), .Y(
        N1285) );
  AOI22X1TF U787 ( .A0(N311), .A1(N1379), .B0(N269), .B1(N35), .Y(N1284) );
  AOI22X1TF U788 ( .A0(N317), .A1(\GR[0][11] ), .B0(N275), .B1(IO_DATAOUTA[11]), .Y(N1283) );
  AOI22X1TF U789 ( .A0(N349), .A1(\GR[5][11] ), .B0(N427), .B1(\GR[7][11] ), 
        .Y(N1214) );
  AOI22X1TF U790 ( .A0(N232), .A1(N1393), .B0(N282), .B1(\GR[6][11] ), .Y(
        N1213) );
  AOI22X1TF U791 ( .A0(N292), .A1(N1379), .B0(N271), .B1(N35), .Y(N1212) );
  AOI22X1TF U792 ( .A0(N230), .A1(\GR[0][11] ), .B0(N284), .B1(IO_DATAOUTA[11]), .Y(N1211) );
  AOI22X1TF U793 ( .A0(N351), .A1(IO_OFFSET[4]), .B0(N286), .B1(\GR[6][4] ), 
        .Y(N1257) );
  AOI22X1TF U794 ( .A0(N311), .A1(\IO_CONTROL[4] ), .B0(N269), .B1(N30), .Y(
        N1256) );
  AOI22X1TF U795 ( .A0(N317), .A1(\GR[0][4] ), .B0(N275), .B1(N26), .Y(N1255)
         );
  AOI22X1TF U796 ( .A0(N349), .A1(\GR[5][4] ), .B0(N427), .B1(\GR[7][4] ), .Y(
        N1186) );
  AOI22X1TF U797 ( .A0(N232), .A1(IO_OFFSET[4]), .B0(N282), .B1(\GR[6][4] ), 
        .Y(N1185) );
  AOI22X1TF U798 ( .A0(N309), .A1(\IO_CONTROL[4] ), .B0(N271), .B1(N30), .Y(
        N1184) );
  AOI22X1TF U799 ( .A0(N230), .A1(\GR[0][4] ), .B0(N284), .B1(N26), .Y(N1183)
         );
  AOI22X1TF U800 ( .A0(N351), .A1(IO_OFFSET[2]), .B0(N285), .B1(\GR[6][2] ), 
        .Y(N1249) );
  AOI22X1TF U801 ( .A0(N349), .A1(\GR[5][2] ), .B0(N427), .B1(\GR[7][2] ), .Y(
        N1178) );
  AOI22X1TF U802 ( .A0(N351), .A1(IO_OFFSET[7]), .B0(N286), .B1(\GR[6][7] ), 
        .Y(N1269) );
  AOI22X1TF U803 ( .A0(N311), .A1(\IO_CONTROL[7] ), .B0(N269), .B1(
        IO_DATAOUTB[7]), .Y(N1268) );
  AOI22X1TF U804 ( .A0(N317), .A1(\GR[0][7] ), .B0(N275), .B1(N28), .Y(N1267)
         );
  AOI22X1TF U805 ( .A0(N349), .A1(\GR[5][7] ), .B0(N427), .B1(\GR[7][7] ), .Y(
        N1198) );
  AOI22X1TF U806 ( .A0(N232), .A1(IO_OFFSET[7]), .B0(N282), .B1(\GR[6][7] ), 
        .Y(N1197) );
  AOI22X1TF U807 ( .A0(N309), .A1(\IO_CONTROL[7] ), .B0(N271), .B1(
        IO_DATAOUTB[7]), .Y(N1196) );
  AOI22X1TF U808 ( .A0(N230), .A1(\GR[0][7] ), .B0(N284), .B1(N28), .Y(N1195)
         );
  AOI22X1TF U809 ( .A0(N351), .A1(IO_OFFSET[8]), .B0(N286), .B1(\GR[6][8] ), 
        .Y(N1273) );
  AOI22X1TF U810 ( .A0(N311), .A1(N1382), .B0(N269), .B1(IO_DATAOUTB[8]), .Y(
        N1272) );
  AOI22X1TF U811 ( .A0(N317), .A1(\GR[0][8] ), .B0(N275), .B1(N31), .Y(N1271)
         );
  AOI22X1TF U812 ( .A0(N349), .A1(\GR[5][8] ), .B0(N1165), .B1(\GR[7][8] ), 
        .Y(N1202) );
  AOI22X1TF U813 ( .A0(N232), .A1(IO_OFFSET[8]), .B0(N281), .B1(\GR[6][8] ), 
        .Y(N1201) );
  AOI22X1TF U814 ( .A0(N309), .A1(N1382), .B0(N270), .B1(IO_DATAOUTB[8]), .Y(
        N1200) );
  AOI22X1TF U815 ( .A0(N230), .A1(\GR[0][8] ), .B0(N283), .B1(N31), .Y(N1199)
         );
  AOI22X1TF U816 ( .A0(N1234), .A1(IO_OFFSET[6]), .B0(N285), .B1(\GR[6][6] ), 
        .Y(N1265) );
  AOI22X1TF U817 ( .A0(N316), .A1(\GR[0][6] ), .B0(N274), .B1(N27), .Y(N1263)
         );
  AOI22X1TF U818 ( .A0(N349), .A1(\GR[5][6] ), .B0(N427), .B1(\GR[7][6] ), .Y(
        N1194) );
  AOI22X1TF U819 ( .A0(N351), .A1(N1394), .B0(N286), .B1(\GR[6][10] ), .Y(
        N1281) );
  AOI22X1TF U820 ( .A0(N311), .A1(N1380), .B0(N269), .B1(IO_DATAOUTB[10]), .Y(
        N1280) );
  AOI22X1TF U821 ( .A0(N317), .A1(\GR[0][10] ), .B0(N275), .B1(N33), .Y(N1279)
         );
  AOI22X1TF U822 ( .A0(N349), .A1(\GR[5][10] ), .B0(N427), .B1(\GR[7][10] ), 
        .Y(N1210) );
  AOI22X1TF U823 ( .A0(N231), .A1(N1394), .B0(N281), .B1(\GR[6][10] ), .Y(
        N1209) );
  AOI22X1TF U824 ( .A0(N309), .A1(N1380), .B0(N270), .B1(IO_DATAOUTB[10]), .Y(
        N1208) );
  AOI22X1TF U825 ( .A0(N229), .A1(\GR[0][10] ), .B0(N283), .B1(N33), .Y(N1207)
         );
  AOI22X1TF U826 ( .A0(N310), .A1(\IO_CONTROL[0] ), .B0(N268), .B1(
        IO_DATAOUTB[0]), .Y(N1240) );
  AOI22X1TF U827 ( .A0(N316), .A1(\GR[0][0] ), .B0(N274), .B1(IO_DATAOUTA[0]), 
        .Y(N1239) );
  AOI22X1TF U828 ( .A0(N1164), .A1(\GR[5][0] ), .B0(N427), .B1(\GR[7][0] ), 
        .Y(N1170) );
  AOI22X1TF U829 ( .A0(N292), .A1(\IO_CONTROL[0] ), .B0(N270), .B1(
        IO_DATAOUTB[0]), .Y(N1168) );
  AOI22X1TF U830 ( .A0(N1148), .A1(N92), .B0(N225), .B1(N250), .Y(N1146) );
  AOI22X1TF U831 ( .A0(N312), .A1(N1378), .B0(N272), .B1(IO_DATAOUTB[12]), .Y(
        N1360) );
  AOI22X1TF U832 ( .A0(N314), .A1(\GR[0][12] ), .B0(N276), .B1(N34), .Y(N1359)
         );
  AOI22X1TF U833 ( .A0(N1148), .A1(N97), .B0(N225), .B1(N252), .Y(N1144) );
  AOI22X1TF U834 ( .A0(N312), .A1(N1380), .B0(N272), .B1(IO_DATAOUTB[10]), .Y(
        N1352) );
  AOI22X1TF U835 ( .A0(N314), .A1(\GR[0][10] ), .B0(N276), .B1(N33), .Y(N1351)
         );
  AOI22X1TF U836 ( .A0(N1148), .A1(N95), .B0(N224), .B1(N254), .Y(N1142) );
  AOI22X1TF U837 ( .A0(N312), .A1(N1382), .B0(N272), .B1(IO_DATAOUTB[8]), .Y(
        N1344) );
  AOI22X1TF U838 ( .A0(N314), .A1(\GR[0][8] ), .B0(N276), .B1(N31), .Y(N1343)
         );
  AOI22X1TF U839 ( .A0(N1148), .A1(N94), .B0(N224), .B1(N248), .Y(N1149) );
  AOI22X1TF U840 ( .A0(N312), .A1(N1376), .B0(N272), .B1(N1387), .Y(N1368) );
  AOI22X1TF U841 ( .A0(N314), .A1(\GR[0][14] ), .B0(N276), .B1(N1384), .Y(
        N1367) );
  AOI22X1TF U842 ( .A0(N1148), .A1(N96), .B0(N225), .B1(N253), .Y(N1143) );
  AOI22X1TF U843 ( .A0(N312), .A1(N1381), .B0(N272), .B1(IO_DATAOUTB[9]), .Y(
        N1348) );
  AOI22X1TF U844 ( .A0(N314), .A1(\GR[0][9] ), .B0(N276), .B1(N32), .Y(N1347)
         );
  AOI22X1TF U845 ( .A0(N1148), .A1(N93), .B0(N225), .B1(N249), .Y(N1147) );
  AOI22X1TF U846 ( .A0(N312), .A1(N1377), .B0(N272), .B1(N1388), .Y(N1364) );
  AOI22X1TF U847 ( .A0(N314), .A1(\GR[0][13] ), .B0(N276), .B1(N1385), .Y(
        N1363) );
  AOI22X1TF U848 ( .A0(N1306), .A1(IO_OFFSET[7]), .B0(N291), .B1(\GR[6][7] ), 
        .Y(N1341) );
  AOI22X1TF U849 ( .A0(N313), .A1(\IO_CONTROL[7] ), .B0(N273), .B1(
        IO_DATAOUTB[7]), .Y(N1340) );
  AOI22X1TF U850 ( .A0(N315), .A1(\GR[0][7] ), .B0(N277), .B1(N28), .Y(N1339)
         );
  AOI22X1TF U851 ( .A0(N224), .A1(N262), .B0(N95), .B1(N1133), .Y(N1130) );
  AOI22X1TF U852 ( .A0(N1306), .A1(IO_OFFSET[0]), .B0(N290), .B1(\GR[6][0] ), 
        .Y(N1313) );
  AOI22X1TF U853 ( .A0(N313), .A1(\IO_CONTROL[0] ), .B0(N273), .B1(
        IO_DATAOUTB[0]), .Y(N1312) );
  AOI22X1TF U854 ( .A0(N314), .A1(\GR[0][0] ), .B0(N276), .B1(IO_DATAOUTA[0]), 
        .Y(N1311) );
  AOI22X1TF U855 ( .A0(N224), .A1(N260), .B0(N97), .B1(N1133), .Y(N1132) );
  AOI22X1TF U856 ( .A0(N350), .A1(IO_OFFSET[2]), .B0(N291), .B1(\GR[6][2] ), 
        .Y(N1321) );
  AOI22X1TF U857 ( .A0(N224), .A1(N261), .B0(N96), .B1(N1133), .Y(N1131) );
  AOI22X1TF U858 ( .A0(N350), .A1(IO_OFFSET[1]), .B0(N291), .B1(\GR[6][1] ), 
        .Y(N1317) );
  AOI22X1TF U859 ( .A0(N313), .A1(\IO_CONTROL[1] ), .B0(N273), .B1(
        IO_DATAOUTB[1]), .Y(N1316) );
  AOI22X1TF U860 ( .A0(N315), .A1(\GR[0][1] ), .B0(N277), .B1(N24), .Y(N1315)
         );
  AOI22X1TF U861 ( .A0(N350), .A1(IO_OFFSET[3]), .B0(N291), .B1(\GR[6][3] ), 
        .Y(N1325) );
  AOI22X1TF U862 ( .A0(N313), .A1(\IO_CONTROL[3] ), .B0(N273), .B1(N29), .Y(
        N1324) );
  AOI22X1TF U863 ( .A0(N315), .A1(\GR[0][3] ), .B0(N277), .B1(IO_DATAOUTA[3]), 
        .Y(N1323) );
  AOI22X1TF U864 ( .A0(N2130), .A1(N1031), .B0(N616), .B1(N977), .Y(N978) );
  AOI22X1TF U865 ( .A0(N2130), .A1(N828), .B0(N330), .B1(N966), .Y(N829) );
  AOI22X1TF U866 ( .A0(N2140), .A1(N1011), .B0(N616), .B1(N1010), .Y(N1012) );
  AOI21X1TF U867 ( .A0(N2220), .A1(N616), .B0(N201), .Y(N984) );
  OAI21X1TF U868 ( .A0(N771), .A1(N542), .B0(N2140), .Y(N543) );
  INVX2TF U869 ( .A(N1122), .Y(N1094) );
  AOI32XLTF U870 ( .A0(N546), .A1(N409), .A2(STATE[3]), .B0(N644), .B1(N545), 
        .Y(N645) );
  AOI21XLTF U871 ( .A0(N752), .A1(N653), .B0(STATE[1]), .Y(N644) );
  OAI32XLTF U872 ( .A0(N22), .A1(CODE_TYPE[1]), .A2(N390), .B0(N1129), .B1(N22), .Y(N1117) );
  MXI2X1TF U873 ( .A(N592), .B(N416), .S0(N1040), .Y(N288) );
  AOI32XLTF U874 ( .A0(CF), .A1(CODE_TYPE[2]), .A2(N372), .B0(N377), .B1(
        CODE_TYPE[2]), .Y(N651) );
  AOI211XLTF U875 ( .A0(N409), .A1(N752), .B0(N546), .C0(N395), .Y(N658) );
  OAI2BB1X1TF U876 ( .A0N(N279), .A1N(N502), .B0(N514), .Y(N1036) );
  OAI2BB1X1TF U877 ( .A0N(N464), .A1N(N580), .B0(N982), .Y(N554) );
  AO21X1TF U878 ( .A0(N615), .A1(N579), .B0(N5750), .Y(N582) );
  OAI2BB1X1TF U879 ( .A0N(N425), .A1N(N465), .B0(N964), .Y(N537) );
  OAI2BB1X1TF U880 ( .A0N(N279), .A1N(N500), .B0(N510), .Y(N1019) );
  OAI2BB1X1TF U881 ( .A0N(N495), .A1N(N279), .B0(N533), .Y(N534) );
  NAND3BX1TF U882 ( .AN(N794), .B(N531), .C(N530), .Y(N1072) );
  NAND2X1TF U883 ( .A(N1018), .B(N786), .Y(N530) );
  OAI2BB2XLTF U884 ( .B0(N1024), .B1(N796), .A0N(N459), .A1N(N425), .Y(N529)
         );
  OAI2BB1X1TF U885 ( .A0N(N494), .A1N(N280), .B0(N556), .Y(N557) );
  OAI222X1TF U886 ( .A0(N199), .A1(N592), .B0(N1078), .B1(N602), .C0(N2560), 
        .C1(N607), .Y(N448) );
  NAND2X1TF U887 ( .A(N471), .B(N580), .Y(N4630) );
  NAND2X1TF U888 ( .A(N595), .B(IO_STATUS[0]), .Y(N587) );
  NOR2BX1TF U889 ( .AN(N584), .B(N1044), .Y(N595) );
  AO22X1TF U890 ( .A0(N562), .A1(REG_A[0]), .B0(N457), .B1(N580), .Y(N563) );
  NAND2X1TF U891 ( .A(N610), .B(REG_A[0]), .Y(N559) );
  XOR2X1TF U892 ( .A(N605), .B(N1064), .Y(N585) );
  OAI2BB1X1TF U893 ( .A0N(REG_B[10]), .A1N(N525), .B0(N524), .Y(N526) );
  OAI2BB1X1TF U894 ( .A0N(N604), .A1N(N1009), .B0(N522), .Y(N523) );
  NAND2BX1TF U895 ( .AN(N1015), .B(N521), .Y(N525) );
  AOI2BB2X1TF U896 ( .B0(N433), .B1(N411), .A0N(N983), .A1N(N411), .Y(N521) );
  NAND2X1TF U897 ( .A(N501), .B(N279), .Y(N528) );
  NAND4X1TF U898 ( .A(N446), .B(N445), .C(N444), .D(N443), .Y(N447) );
  NAND2X1TF U899 ( .A(N618), .B(N2140), .Y(N443) );
  NAND2X1TF U900 ( .A(N965), .B(N616), .Y(N444) );
  AOI2BB2X1TF U901 ( .B0(N442), .B1(REG_A[12]), .A0N(N622), .A1N(N568), .Y(
        N445) );
  AO21X1TF U902 ( .A0(N434), .A1(N568), .B0(N643), .Y(N442) );
  NAND2BX1TF U903 ( .AN(N621), .B(N609), .Y(N446) );
  NAND2X1TF U904 ( .A(N503), .B(N279), .Y(N450) );
  OAI2BB1X1TF U905 ( .A0N(N425), .A1N(N470), .B0(N456), .Y(N4570) );
  OAI2BB2XLTF U906 ( .B0(N454), .B1(N608), .A0N(N604), .A1N(N1011), .Y(N455)
         );
  CLKBUFX2TF U907 ( .A(N373), .Y(N436) );
  NAND3X1TF U908 ( .A(N613), .B(N377), .C(N390), .Y(N648) );
  NAND2X1TF U909 ( .A(CODE_TYPE[1]), .B(N1122), .Y(N1086) );
  NAND3X1TF U910 ( .A(N451), .B(N1085), .C(N614), .Y(N441) );
  INVX2TF U911 ( .A(N623), .Y(N667) );
  NAND2X1TF U912 ( .A(N623), .B(CODE_TYPE[2]), .Y(N451) );
  AO22X1TF U913 ( .A0(N1018), .A1(N1017), .B0(REG_A[9]), .B1(N1016), .Y(N385)
         );
  CLKBUFX2TF U914 ( .A(N1165), .Y(N427) );
  CLKBUFX2TF U915 ( .A(N1237), .Y(N430) );
  CLKBUFX2TF U916 ( .A(N1309), .Y(N432) );
  NAND2X1TF U917 ( .A(REG_A[11]), .B(N641), .Y(N763) );
  NAND2X1TF U918 ( .A(N426), .B(REG_A[10]), .Y(N814) );
  NAND2X1TF U919 ( .A(REG_A[13]), .B(N641), .Y(N632) );
  NAND2X1TF U920 ( .A(N2100), .B(N667), .Y(N1085) );
  NAND3X1TF U921 ( .A(N560), .B(N377), .C(N390), .Y(N1087) );
  NAND2X1TF U922 ( .A(N641), .B(REG_A[7]), .Y(N764) );
  NAND2X1TF U923 ( .A(N807), .B(REG_A[5]), .Y(N783) );
  NAND2X1TF U924 ( .A(N2210), .B(REG_A[8]), .Y(N813) );
  NAND2X1TF U925 ( .A(REG_A[6]), .B(N426), .Y(N819) );
  NAND4X1TF U926 ( .A(N764), .B(N783), .C(N813), .D(N819), .Y(N828) );
  NAND2X1TF U927 ( .A(N641), .B(REG_A[3]), .Y(N784) );
  AOI222XLTF U928 ( .A0(N828), .A1(N988), .B0(N987), .B1(N818), .C0(N963), 
        .C1(N986), .Y(N621) );
  NAND2X1TF U929 ( .A(N426), .B(REG_A[7]), .Y(N772) );
  NAND2X1TF U930 ( .A(N2210), .B(REG_A[9]), .Y(N769) );
  NAND2X1TF U931 ( .A(N333), .B(REG_A[8]), .Y(N800) );
  NAND2X1TF U932 ( .A(REG_A[6]), .B(N807), .Y(N624) );
  NAND4X1TF U933 ( .A(N772), .B(N769), .C(N800), .D(N624), .Y(N1011) );
  NAND2X1TF U934 ( .A(N641), .B(REG_A[4]), .Y(N798) );
  OAI221XLTF U935 ( .A0(N371), .A1(REG_A[0]), .B0(REG_B[0]), .B1(REG_A[1]), 
        .C0(N406), .Y(N994) );
  AOI2BB2X1TF U936 ( .B0(N1021), .B1(N197), .A0N(N197), .A1N(N994), .Y(N779)
         );
  NAND2X1TF U937 ( .A(REG_B[3]), .B(N609), .Y(N627) );
  OAI222X1TF U938 ( .A0(N1078), .A1(N605), .B0(N199), .B1(N6030), .C0(N2600), 
        .C1(N607), .Y(N368) );
  NAND2X1TF U939 ( .A(REG_A[12]), .B(N343), .Y(N633) );
  NAND2X1TF U940 ( .A(N789), .B(N197), .Y(N768) );
  NAND2X1TF U941 ( .A(N407), .B(N790), .Y(N1004) );
  NAND2X1TF U942 ( .A(N426), .B(REG_A[8]), .Y(N765) );
  NAND2X1TF U943 ( .A(N807), .B(REG_A[7]), .Y(N821) );
  NAND2X1TF U944 ( .A(N641), .B(REG_A[9]), .Y(N815) );
  NAND4X1TF U945 ( .A(N635), .B(N765), .C(N821), .D(N815), .Y(N1006) );
  NAND2X1TF U946 ( .A(N641), .B(REG_A[5]), .Y(N822) );
  NAND2X1TF U947 ( .A(REG_A[6]), .B(N2210), .Y(N767) );
  AOI222XLTF U948 ( .A0(N1006), .A1(N988), .B0(N787), .B1(N987), .C0(N1009), 
        .C1(N986), .Y(N637) );
  OAI222X1TF U949 ( .A0(N1078), .A1(N6030), .B0(N199), .B1(N602), .C0(N2570), 
        .C1(N607), .Y(N438) );
  NAND2X1TF U950 ( .A(N807), .B(REG_A[8]), .Y(N773) );
  NAND2X1TF U951 ( .A(N641), .B(REG_A[10]), .Y(N770) );
  NAND2X1TF U952 ( .A(N343), .B(REG_A[9]), .Y(N801) );
  NAND4X1TF U953 ( .A(N773), .B(N770), .C(N801), .D(N639), .Y(N1023) );
  NAND2X1TF U954 ( .A(REG_A[6]), .B(N641), .Y(N774) );
  NAND2X1TF U955 ( .A(N2220), .B(REG_A[7]), .Y(N802) );
  NAND2X1TF U956 ( .A(N343), .B(REG_A[5]), .Y(N797) );
  NAND2X1TF U957 ( .A(N807), .B(REG_A[4]), .Y(N640) );
  NAND4X1TF U958 ( .A(N774), .B(N802), .C(N797), .D(N640), .Y(N1031) );
  NAND2X1TF U959 ( .A(N333), .B(REG_A[2]), .Y(N991) );
  NAND2X1TF U960 ( .A(N370), .B(N752), .Y(N754) );
  NAND2X1TF U961 ( .A(N546), .B(START), .Y(N653) );
  NOR2BX1TF U962 ( .AN(N758), .B(N690), .Y(N166) );
  NAND2X1TF U963 ( .A(I_ADDR[1]), .B(I_ADDR[2]), .Y(N727) );
  NAND2X1TF U964 ( .A(N730), .B(I_ADDR[4]), .Y(N733) );
  NAND2X1TF U965 ( .A(N736), .B(I_ADDR[6]), .Y(N739) );
  NAND2X1TF U966 ( .A(N743), .B(I_ADDR[8]), .Y(N742) );
  AO22X1TF U967 ( .A0(I_ADDR[0]), .A1(SMDR[8]), .B0(N412), .B1(SMDR[0]), .Y(
        D_DATAOUT[0]) );
  AO22X1TF U968 ( .A0(I_ADDR[0]), .A1(SMDR[9]), .B0(N412), .B1(SMDR[1]), .Y(
        D_DATAOUT[1]) );
  AO22X1TF U969 ( .A0(I_ADDR[0]), .A1(SMDR[10]), .B0(N412), .B1(SMDR[2]), .Y(
        D_DATAOUT[2]) );
  AO22X1TF U970 ( .A0(I_ADDR[0]), .A1(SMDR[11]), .B0(N412), .B1(SMDR[3]), .Y(
        D_DATAOUT[3]) );
  AO22X1TF U971 ( .A0(I_ADDR[0]), .A1(SMDR[12]), .B0(N412), .B1(SMDR[4]), .Y(
        D_DATAOUT[4]) );
  AO22X1TF U972 ( .A0(I_ADDR[0]), .A1(SMDR[13]), .B0(N412), .B1(SMDR[5]), .Y(
        D_DATAOUT[5]) );
  AO22X1TF U973 ( .A0(I_ADDR[0]), .A1(SMDR[14]), .B0(N412), .B1(SMDR[6]), .Y(
        D_DATAOUT[6]) );
  AO22X1TF U974 ( .A0(I_ADDR[0]), .A1(SMDR[15]), .B0(N412), .B1(SMDR[7]), .Y(
        D_DATAOUT[7]) );
  NOR4XLTF U975 ( .A(N757), .B(N1124), .C(N658), .D(N412), .Y(N660) );
  OAI221XLTF U976 ( .A0(CODE_TYPE[1]), .A1(N612), .B0(N377), .B1(N384), .C0(
        N560), .Y(N664) );
  AOI2BB2X1TF U977 ( .B0(N246), .B1(N681), .A0N(\GR[0][0] ), .A1N(N245), .Y(
        N958) );
  AOI2BB2X1TF U978 ( .B0(N246), .B1(N682), .A0N(\GR[0][1] ), .A1N(N245), .Y(
        N957) );
  AOI2BB2X1TF U979 ( .B0(N246), .B1(N683), .A0N(\GR[0][2] ), .A1N(N245), .Y(
        N956) );
  AOI2BB2X1TF U980 ( .B0(N246), .B1(N684), .A0N(\GR[0][3] ), .A1N(N245), .Y(
        N955) );
  AOI2BB2X1TF U981 ( .B0(N246), .B1(N685), .A0N(\GR[0][4] ), .A1N(N245), .Y(
        N954) );
  AOI2BB2X1TF U982 ( .B0(N246), .B1(N686), .A0N(\GR[0][5] ), .A1N(N245), .Y(
        N953) );
  AOI2BB2X1TF U983 ( .B0(N246), .B1(N687), .A0N(\GR[0][6] ), .A1N(N245), .Y(
        N952) );
  AOI2BB2X1TF U984 ( .B0(N246), .B1(N688), .A0N(\GR[0][7] ), .A1N(N245), .Y(
        N951) );
  AOI2BB2X1TF U985 ( .B0(N339), .B1(N681), .A0N(\IO_CONTROL[0] ), .A1N(N673), 
        .Y(N950) );
  AOI2BB2X1TF U986 ( .B0(N339), .B1(N682), .A0N(\IO_CONTROL[1] ), .A1N(N673), 
        .Y(N949) );
  AOI2BB2X1TF U987 ( .B0(N339), .B1(N683), .A0N(\IO_CONTROL[2] ), .A1N(N673), 
        .Y(N948) );
  AOI2BB2X1TF U988 ( .B0(N339), .B1(N684), .A0N(\IO_CONTROL[3] ), .A1N(N673), 
        .Y(N947) );
  AOI2BB2X1TF U989 ( .B0(N339), .B1(N685), .A0N(\IO_CONTROL[4] ), .A1N(N673), 
        .Y(N946) );
  AOI2BB2X1TF U990 ( .B0(N339), .B1(N686), .A0N(\IO_CONTROL[5] ), .A1N(N673), 
        .Y(N945) );
  AOI2BB2X1TF U991 ( .B0(N339), .B1(N687), .A0N(\IO_CONTROL[6] ), .A1N(N673), 
        .Y(N944) );
  AOI2BB2X1TF U992 ( .B0(N339), .B1(N688), .A0N(\IO_CONTROL[7] ), .A1N(N673), 
        .Y(N943) );
  AOI2BB2X1TF U993 ( .B0(N340), .B1(N681), .A0N(IO_DATAOUTA[0]), .A1N(N674), 
        .Y(N942) );
  AOI2BB2X1TF U994 ( .B0(N340), .B1(N682), .A0N(N24), .A1N(N674), .Y(N941) );
  AOI2BB2X1TF U995 ( .B0(N340), .B1(N683), .A0N(N25), .A1N(N674), .Y(N940) );
  AOI2BB2X1TF U996 ( .B0(N340), .B1(N684), .A0N(IO_DATAOUTA[3]), .A1N(N674), 
        .Y(N939) );
  AOI2BB2X1TF U997 ( .B0(N340), .B1(N685), .A0N(N26), .A1N(N674), .Y(N938) );
  AOI2BB2X1TF U998 ( .B0(N340), .B1(N686), .A0N(IO_DATAOUTA[5]), .A1N(N674), 
        .Y(N937) );
  AOI2BB2X1TF U999 ( .B0(N340), .B1(N687), .A0N(N27), .A1N(N674), .Y(N936) );
  AOI2BB2X1TF U1000 ( .B0(N340), .B1(N688), .A0N(N28), .A1N(N674), .Y(N935) );
  AOI2BB2X1TF U1001 ( .B0(N267), .B1(N681), .A0N(IO_DATAOUTB[0]), .A1N(N266), 
        .Y(N934) );
  AOI2BB2X1TF U1002 ( .B0(N267), .B1(N682), .A0N(IO_DATAOUTB[1]), .A1N(N266), 
        .Y(N933) );
  AOI2BB2X1TF U1003 ( .B0(N267), .B1(N683), .A0N(IO_DATAOUTB[2]), .A1N(N266), 
        .Y(N932) );
  AOI2BB2X1TF U1004 ( .B0(N267), .B1(N684), .A0N(N29), .A1N(N266), .Y(N931) );
  AOI2BB2X1TF U1005 ( .B0(N267), .B1(N685), .A0N(N30), .A1N(N266), .Y(N930) );
  AOI2BB2X1TF U1006 ( .B0(N267), .B1(N686), .A0N(IO_DATAOUTB[5]), .A1N(N266), 
        .Y(N929) );
  AOI2BB2X1TF U1007 ( .B0(N267), .B1(N687), .A0N(N23), .A1N(N266), .Y(N928) );
  AOI2BB2X1TF U1008 ( .B0(N267), .B1(N688), .A0N(IO_DATAOUTB[7]), .A1N(N266), 
        .Y(N927) );
  AOI2BB2X1TF U1009 ( .B0(N244), .B1(N681), .A0N(IO_OFFSET[0]), .A1N(N243), 
        .Y(N926) );
  AOI2BB2X1TF U1010 ( .B0(N244), .B1(N682), .A0N(IO_OFFSET[1]), .A1N(N243), 
        .Y(N925) );
  AOI2BB2X1TF U1011 ( .B0(N244), .B1(N683), .A0N(IO_OFFSET[2]), .A1N(N243), 
        .Y(N924) );
  AOI2BB2X1TF U1012 ( .B0(N244), .B1(N684), .A0N(IO_OFFSET[3]), .A1N(N243), 
        .Y(N923) );
  AOI2BB2X1TF U1013 ( .B0(N244), .B1(N685), .A0N(IO_OFFSET[4]), .A1N(N243), 
        .Y(N922) );
  AOI2BB2X1TF U1014 ( .B0(N244), .B1(N686), .A0N(IO_OFFSET[5]), .A1N(N243), 
        .Y(N921) );
  AOI2BB2X1TF U1015 ( .B0(N244), .B1(N687), .A0N(IO_OFFSET[6]), .A1N(N243), 
        .Y(N920) );
  AOI2BB2X1TF U1016 ( .B0(N244), .B1(N688), .A0N(IO_OFFSET[7]), .A1N(N243), 
        .Y(N919) );
  AOI2BB2X1TF U1017 ( .B0(N2480), .B1(N681), .A0N(\GR[5][0] ), .A1N(N2470), 
        .Y(N918) );
  AOI2BB2X1TF U1018 ( .B0(N2480), .B1(N682), .A0N(\GR[5][1] ), .A1N(N2470), 
        .Y(N917) );
  AOI2BB2X1TF U1019 ( .B0(N2480), .B1(N683), .A0N(\GR[5][2] ), .A1N(N2470), 
        .Y(N916) );
  AOI2BB2X1TF U1020 ( .B0(N2480), .B1(N684), .A0N(\GR[5][3] ), .A1N(N2470), 
        .Y(N915) );
  AOI2BB2X1TF U1021 ( .B0(N2480), .B1(N685), .A0N(\GR[5][4] ), .A1N(N2470), 
        .Y(N914) );
  AOI2BB2X1TF U1022 ( .B0(N2480), .B1(N686), .A0N(\GR[5][5] ), .A1N(N2470), 
        .Y(N913) );
  AOI2BB2X1TF U1023 ( .B0(N2480), .B1(N687), .A0N(\GR[5][6] ), .A1N(N2470), 
        .Y(N912) );
  AOI2BB2X1TF U1024 ( .B0(N2480), .B1(N688), .A0N(\GR[5][7] ), .A1N(N2470), 
        .Y(N911) );
  AOI2BB2X1TF U1025 ( .B0(N242), .B1(N681), .A0N(\GR[6][0] ), .A1N(N241), .Y(
        N910) );
  AOI2BB2X1TF U1026 ( .B0(N242), .B1(N682), .A0N(\GR[6][1] ), .A1N(N241), .Y(
        N909) );
  AOI2BB2X1TF U1027 ( .B0(N242), .B1(N683), .A0N(\GR[6][2] ), .A1N(N241), .Y(
        N908) );
  AOI2BB2X1TF U1028 ( .B0(N242), .B1(N684), .A0N(\GR[6][3] ), .A1N(N241), .Y(
        N907) );
  AOI2BB2X1TF U1029 ( .B0(N242), .B1(N685), .A0N(\GR[6][4] ), .A1N(N241), .Y(
        N906) );
  AOI2BB2X1TF U1030 ( .B0(N242), .B1(N686), .A0N(\GR[6][5] ), .A1N(N241), .Y(
        N905) );
  AOI2BB2X1TF U1031 ( .B0(N242), .B1(N687), .A0N(\GR[6][6] ), .A1N(N241), .Y(
        N904) );
  AOI2BB2X1TF U1032 ( .B0(N242), .B1(N688), .A0N(\GR[6][7] ), .A1N(N241), .Y(
        N903) );
  AOI2BB2X1TF U1033 ( .B0(N240), .B1(N681), .A0N(\GR[7][0] ), .A1N(N239), .Y(
        N902) );
  AOI2BB2X1TF U1034 ( .B0(N240), .B1(N682), .A0N(\GR[7][1] ), .A1N(N239), .Y(
        N901) );
  AOI2BB2X1TF U1035 ( .B0(N240), .B1(N683), .A0N(\GR[7][2] ), .A1N(N239), .Y(
        N900) );
  AOI2BB2X1TF U1036 ( .B0(N240), .B1(N684), .A0N(\GR[7][3] ), .A1N(N239), .Y(
        N899) );
  AOI2BB2X1TF U1037 ( .B0(N240), .B1(N685), .A0N(\GR[7][4] ), .A1N(N239), .Y(
        N898) );
  AOI2BB2X1TF U1038 ( .B0(N240), .B1(N686), .A0N(\GR[7][5] ), .A1N(N239), .Y(
        N897) );
  AOI2BB2X1TF U1039 ( .B0(N240), .B1(N687), .A0N(\GR[7][6] ), .A1N(N239), .Y(
        N896) );
  AOI2BB2X1TF U1040 ( .B0(N240), .B1(N688), .A0N(\GR[7][7] ), .A1N(N239), .Y(
        N895) );
  AOI2BB2X1TF U1041 ( .B0(N238), .B1(N709), .A0N(\GR[0][8] ), .A1N(N237), .Y(
        N894) );
  AOI2BB2X1TF U1042 ( .B0(N238), .B1(N710), .A0N(\GR[0][9] ), .A1N(N237), .Y(
        N893) );
  AOI2BB2X1TF U1043 ( .B0(N238), .B1(N711), .A0N(\GR[0][10] ), .A1N(N237), .Y(
        N892) );
  AOI2BB2X1TF U1044 ( .B0(N238), .B1(N712), .A0N(\GR[0][11] ), .A1N(N237), .Y(
        N891) );
  AOI2BB2X1TF U1045 ( .B0(N238), .B1(N714), .A0N(\GR[0][12] ), .A1N(N237), .Y(
        N890) );
  AOI2BB2X1TF U1046 ( .B0(N238), .B1(N715), .A0N(\GR[0][13] ), .A1N(N237), .Y(
        N889) );
  AOI2BB2X1TF U1047 ( .B0(N238), .B1(N716), .A0N(\GR[0][14] ), .A1N(N237), .Y(
        N888) );
  AOI2BB2X1TF U1048 ( .B0(N238), .B1(N723), .A0N(\GR[0][15] ), .A1N(N237), .Y(
        N887) );
  AOI2BB2X1TF U1049 ( .B0(N263), .B1(N709), .A0N(N1382), .A1N(N2530), .Y(N886)
         );
  AOI2BB2X1TF U1050 ( .B0(N263), .B1(N710), .A0N(N1381), .A1N(N2530), .Y(N885)
         );
  AOI2BB2X1TF U1051 ( .B0(N263), .B1(N711), .A0N(N1380), .A1N(N2530), .Y(N884)
         );
  AOI2BB2X1TF U1052 ( .B0(N263), .B1(N712), .A0N(N1379), .A1N(N2530), .Y(N883)
         );
  AOI2BB2X1TF U1053 ( .B0(N263), .B1(N714), .A0N(N1378), .A1N(N2530), .Y(N8820) );
  AOI2BB2X1TF U1054 ( .B0(N263), .B1(N715), .A0N(N1377), .A1N(N2530), .Y(N881)
         );
  AOI2BB2X1TF U1055 ( .B0(N263), .B1(N716), .A0N(N1376), .A1N(N2530), .Y(N880)
         );
  AOI2BB2X1TF U1056 ( .B0(N263), .B1(N723), .A0N(N1375), .A1N(N2530), .Y(N879)
         );
  AOI2BB2X1TF U1057 ( .B0(N265), .B1(N709), .A0N(N31), .A1N(N264), .Y(N878) );
  AOI2BB2X1TF U1058 ( .B0(N265), .B1(N710), .A0N(N32), .A1N(N265), .Y(N877) );
  AOI2BB2X1TF U1059 ( .B0(N265), .B1(N711), .A0N(N33), .A1N(N264), .Y(N876) );
  AOI2BB2X1TF U1060 ( .B0(N265), .B1(N712), .A0N(IO_DATAOUTA[11]), .A1N(N264), 
        .Y(N875) );
  AOI2BB2X1TF U1061 ( .B0(N265), .B1(N714), .A0N(N34), .A1N(N264), .Y(N874) );
  AOI2BB2X1TF U1062 ( .B0(N265), .B1(N715), .A0N(N1385), .A1N(N264), .Y(N873)
         );
  AOI2BB2X1TF U1063 ( .B0(N265), .B1(N716), .A0N(N1384), .A1N(N264), .Y(N872)
         );
  AOI2BB2X1TF U1064 ( .B0(N264), .B1(N723), .A0N(N1383), .A1N(N264), .Y(N871)
         );
  AOI2BB2X1TF U1065 ( .B0(N2500), .B1(N709), .A0N(IO_DATAOUTB[8]), .A1N(N2490), 
        .Y(N870) );
  AOI2BB2X1TF U1066 ( .B0(N2500), .B1(N710), .A0N(IO_DATAOUTB[9]), .A1N(N2490), 
        .Y(N869) );
  AOI2BB2X1TF U1067 ( .B0(N2500), .B1(N711), .A0N(IO_DATAOUTB[10]), .A1N(N2490), .Y(N868) );
  AOI2BB2X1TF U1068 ( .B0(N2500), .B1(N712), .A0N(N35), .A1N(N2490), .Y(N867)
         );
  AOI2BB2X1TF U1069 ( .B0(N2500), .B1(N714), .A0N(IO_DATAOUTB[12]), .A1N(N2490), .Y(N866) );
  AOI2BB2X1TF U1070 ( .B0(N2500), .B1(N715), .A0N(N1388), .A1N(N2490), .Y(N865) );
  AOI2BB2X1TF U1071 ( .B0(N2500), .B1(N716), .A0N(N1387), .A1N(N2490), .Y(N864) );
  AOI2BB2X1TF U1072 ( .B0(N2500), .B1(N723), .A0N(N1386), .A1N(N2490), .Y(N863) );
  AOI2BB2X1TF U1073 ( .B0(N337), .B1(N709), .A0N(IO_OFFSET[8]), .A1N(N702), 
        .Y(N862) );
  AOI2BB2X1TF U1074 ( .B0(N337), .B1(N710), .A0N(IO_OFFSET[9]), .A1N(N702), 
        .Y(N861) );
  AOI2BB2X1TF U1075 ( .B0(N337), .B1(N711), .A0N(N1394), .A1N(N702), .Y(N860)
         );
  AOI2BB2X1TF U1076 ( .B0(N337), .B1(N712), .A0N(N1393), .A1N(N702), .Y(N859)
         );
  AOI2BB2X1TF U1077 ( .B0(N337), .B1(N714), .A0N(N1392), .A1N(N702), .Y(N858)
         );
  AOI2BB2X1TF U1078 ( .B0(N337), .B1(N715), .A0N(N1391), .A1N(N702), .Y(N857)
         );
  AOI2BB2X1TF U1079 ( .B0(N337), .B1(N716), .A0N(N1390), .A1N(N702), .Y(N856)
         );
  AOI2BB2X1TF U1080 ( .B0(N337), .B1(N723), .A0N(N1389), .A1N(N702), .Y(N855)
         );
  AOI2BB2X1TF U1081 ( .B0(N2520), .B1(N709), .A0N(\GR[5][8] ), .A1N(N2510), 
        .Y(N854) );
  AOI2BB2X1TF U1082 ( .B0(N2520), .B1(N710), .A0N(\GR[5][9] ), .A1N(N2510), 
        .Y(N853) );
  AOI2BB2X1TF U1083 ( .B0(N2520), .B1(N711), .A0N(\GR[5][10] ), .A1N(N2510), 
        .Y(N852) );
  AOI2BB2X1TF U1084 ( .B0(N2520), .B1(N712), .A0N(\GR[5][11] ), .A1N(N2510), 
        .Y(N851) );
  AOI2BB2X1TF U1085 ( .B0(N2520), .B1(N714), .A0N(\GR[5][12] ), .A1N(N2510), 
        .Y(N850) );
  AOI2BB2X1TF U1086 ( .B0(N2520), .B1(N715), .A0N(\GR[5][13] ), .A1N(N2510), 
        .Y(N849) );
  AOI2BB2X1TF U1087 ( .B0(N2520), .B1(N716), .A0N(\GR[5][14] ), .A1N(N2510), 
        .Y(N848) );
  AOI2BB2X1TF U1088 ( .B0(N2520), .B1(N723), .A0N(\GR[5][15] ), .A1N(N2510), 
        .Y(N847) );
  AOI2BB2X1TF U1089 ( .B0(N236), .B1(N709), .A0N(\GR[6][8] ), .A1N(N235), .Y(
        N846) );
  AOI2BB2X1TF U1090 ( .B0(N236), .B1(N710), .A0N(\GR[6][9] ), .A1N(N235), .Y(
        N845) );
  AOI2BB2X1TF U1091 ( .B0(N236), .B1(N711), .A0N(\GR[6][10] ), .A1N(N235), .Y(
        N844) );
  AOI2BB2X1TF U1092 ( .B0(N236), .B1(N712), .A0N(\GR[6][11] ), .A1N(N235), .Y(
        N843) );
  AOI2BB2X1TF U1093 ( .B0(N236), .B1(N714), .A0N(\GR[6][12] ), .A1N(N235), .Y(
        N842) );
  AOI2BB2X1TF U1094 ( .B0(N236), .B1(N715), .A0N(\GR[6][13] ), .A1N(N235), .Y(
        N841) );
  AOI2BB2X1TF U1095 ( .B0(N236), .B1(N716), .A0N(\GR[6][14] ), .A1N(N235), .Y(
        N840) );
  AOI2BB2X1TF U1096 ( .B0(N236), .B1(N723), .A0N(\GR[6][15] ), .A1N(N235), .Y(
        N839) );
  AOI2BB2X1TF U1097 ( .B0(N336), .B1(N709), .A0N(\GR[7][8] ), .A1N(N724), .Y(
        N838) );
  AOI2BB2X1TF U1098 ( .B0(N336), .B1(N710), .A0N(\GR[7][9] ), .A1N(N724), .Y(
        N837) );
  AOI2BB2X1TF U1099 ( .B0(N336), .B1(N711), .A0N(\GR[7][10] ), .A1N(N724), .Y(
        N836) );
  AOI2BB2X1TF U1100 ( .B0(N336), .B1(N712), .A0N(\GR[7][11] ), .A1N(N724), .Y(
        N835) );
  AOI2BB2X1TF U1101 ( .B0(N336), .B1(N714), .A0N(\GR[7][12] ), .A1N(N724), .Y(
        N834) );
  AOI2BB2X1TF U1102 ( .B0(N336), .B1(N715), .A0N(\GR[7][13] ), .A1N(N724), .Y(
        N833) );
  AOI2BB2X1TF U1103 ( .B0(N336), .B1(N716), .A0N(\GR[7][14] ), .A1N(N724), .Y(
        N832) );
  AOI2BB2X1TF U1104 ( .B0(N336), .B1(N723), .A0N(\GR[7][15] ), .A1N(N724), .Y(
        N831) );
  NOR4XLTF U1105 ( .A(\IO_CONTROL[4] ), .B(\IO_CONTROL[5] ), .C(
        \IO_CONTROL[6] ), .D(\IO_CONTROL[7] ), .Y(N753) );
  NOR4XLTF U1106 ( .A(IO_STATUS[0]), .B(IO_STATUS[1]), .C(IO_STATUS[2]), .D(
        N753), .Y(N755) );
  NAND2X1TF U1108 ( .A(N988), .B(N790), .Y(N1028) );
  NAND2X1TF U1109 ( .A(N807), .B(REG_A[9]), .Y(N766) );
  NAND4X1TF U1110 ( .A(N767), .B(N766), .C(N765), .D(N764), .Y(N786) );
  NAND4BX1TF U1111 ( .AN(N777), .B(N774), .C(N773), .D(N772), .Y(N989) );
  OAI2BB2XLTF U1112 ( .B0(N778), .B1(N387), .A0N(N989), .A1N(N616), .Y(N781)
         );
  NAND2X1TF U1113 ( .A(N609), .B(N407), .Y(N995) );
  NAND2X1TF U1114 ( .A(N790), .B(N986), .Y(N979) );
  OA21XLTF U1115 ( .A0(N436), .A1(REG_B[2]), .B0(N984), .Y(N793) );
  NAND4BX1TF U1116 ( .AN(N803), .B(N802), .C(N801), .D(N800), .Y(N977) );
  AOI2BB2X1TF U1117 ( .B0(N1018), .B1(N977), .A0N(N979), .A1N(N1025), .Y(N812)
         );
  NAND2X1TF U1118 ( .A(N2220), .B(REG_A[15]), .Y(N1027) );
  AOI2BB2X1TF U1119 ( .B0(REG_A[3]), .B1(N810), .A0N(N407), .A1N(N809), .Y(
        N811) );
  NAND4BX1TF U1120 ( .AN(N816), .B(N815), .C(N814), .D(N813), .Y(N966) );
  OAI2BB2XLTF U1121 ( .B0(N817), .B1(N393), .A0N(N966), .A1N(N1018), .Y(N825)
         );
  NAND2X1TF U1122 ( .A(N2220), .B(REG_A[4]), .Y(N820) );
  NAND4X1TF U1123 ( .A(N822), .B(N821), .C(N820), .D(N819), .Y(N967) );
  AOI2BB2X1TF U1124 ( .B0(N616), .B1(N967), .A0N(N979), .A1N(N827), .Y(N823)
         );
  NAND2X1TF U1125 ( .A(N609), .B(N986), .Y(N1029) );
  AOI222XLTF U1126 ( .A0(N967), .A1(N988), .B0(N966), .B1(N986), .C0(N965), 
        .C1(N987), .Y(N974) );
  OAI221XLTF U1127 ( .A0(REG_A[1]), .A1(N373), .B0(N386), .B1(N983), .C0(N615), 
        .Y(N1002) );
  AOI222XLTF U1128 ( .A0(N989), .A1(N988), .B0(N1017), .B1(N987), .C0(N1010), 
        .C1(N986), .Y(N999) );
  NAND2X1TF U1129 ( .A(N343), .B(REG_A[3]), .Y(N992) );
  NAND2BX1TF U1130 ( .AN(N994), .B(N197), .Y(N1013) );
  AOI2BB2X1TF U1131 ( .B0(N616), .B1(N996), .A0N(N995), .A1N(N1013), .Y(N997)
         );
  AO21X1TF U1132 ( .A0(N435), .A1(N570), .B0(N200), .Y(N1007) );
  AO21X1TF U1133 ( .A0(N435), .A1(N571), .B0(N201), .Y(N1016) );
  OAI2BB2XLTF U1134 ( .B0(N1025), .B1(N1024), .A0N(N1023), .A1N(N2140), .Y(
        N1038) );
  NAND3X1TF U1135 ( .A(N1047), .B(N1046), .C(N1045), .Y(N328) );
  AOI2BB2X1TF U1136 ( .B0(IO_DATAINA[9]), .B1(N2160), .A0N(N607), .A1N(N2620), 
        .Y(N1052) );
  AOI2BB2X1TF U1137 ( .B0(IO_DATAINA[12]), .B1(N2160), .A0N(N607), .A1N(N2610), 
        .Y(N1055) );
  AOI2BB2X1TF U1138 ( .B0(IO_DATAINA[11]), .B1(N2160), .A0N(N607), .A1N(N2590), 
        .Y(N1062) );
  AOI2BB2X1TF U1139 ( .B0(IO_DATAINA[10]), .B1(N2160), .A0N(N607), .A1N(N2580), 
        .Y(N1066) );
  OAI2BB2XLTF U1140 ( .B0(N22), .B1(N1091), .A0N(N1120), .A1N(N613), .Y(N1092)
         );
  AOI2BB2X1TF U1141 ( .B0(N225), .B1(N255), .A0N(N2550), .A1N(N1140), .Y(N1141) );
  AOI2BB2X1TF U1142 ( .B0(N225), .B1(N251), .A0N(N2540), .A1N(N1150), .Y(N1145) );
  AOI2BB2X1TF U1143 ( .B0(N225), .B1(N247), .A0N(N2550), .A1N(N1150), .Y(N1151) );
  NAND4X1TF U1144 ( .A(N1167), .B(N1168), .C(N1169), .D(N1170), .Y(N185) );
  NAND4X1TF U1145 ( .A(N1171), .B(N1172), .C(N1173), .D(N1174), .Y(N184) );
  NAND4X1TF U1146 ( .A(N1175), .B(N1176), .C(N1177), .D(N1178), .Y(N183) );
  NAND4X1TF U1147 ( .A(N1179), .B(N1180), .C(N1181), .D(N1182), .Y(N182) );
  NAND4X1TF U1148 ( .A(N1183), .B(N1184), .C(N1185), .D(N1186), .Y(N181) );
  NAND4X1TF U1149 ( .A(N1187), .B(N1188), .C(N1189), .D(N1190), .Y(N180) );
  NAND4X1TF U1150 ( .A(N1191), .B(N1192), .C(N1193), .D(N1194), .Y(N179) );
  NAND4X1TF U1151 ( .A(N1195), .B(N1196), .C(N1197), .D(N1198), .Y(N178) );
  NAND4X1TF U1152 ( .A(N1199), .B(N1200), .C(N1201), .D(N1202), .Y(N177) );
  NAND4X1TF U1153 ( .A(N1203), .B(N1204), .C(N1205), .D(N1206), .Y(N176) );
  NAND4X1TF U1154 ( .A(N1207), .B(N1208), .C(N1209), .D(N1210), .Y(N175) );
  NAND4X1TF U1155 ( .A(N1211), .B(N1212), .C(N1213), .D(N1214), .Y(N174) );
  NAND4X1TF U1156 ( .A(N1215), .B(N1216), .C(N1217), .D(N1218), .Y(N173) );
  NAND4X1TF U1157 ( .A(N1219), .B(N1220), .C(N1221), .D(N1222), .Y(N172) );
  NAND4X1TF U1158 ( .A(N1223), .B(N1224), .C(N1225), .D(N1226), .Y(N171) );
  NAND4X1TF U1159 ( .A(N1227), .B(N1228), .C(N1229), .D(N1230), .Y(N170) );
  NAND4X1TF U1160 ( .A(N1239), .B(N1240), .C(N1241), .D(N1242), .Y(N222) );
  NAND4X1TF U1161 ( .A(N1243), .B(N1244), .C(N1245), .D(N1246), .Y(N221) );
  NAND4X1TF U1162 ( .A(N1247), .B(N1248), .C(N1249), .D(N1250), .Y(N220) );
  NAND4X1TF U1163 ( .A(N1251), .B(N1252), .C(N1253), .D(N1254), .Y(N219) );
  NAND4X1TF U1164 ( .A(N1255), .B(N1256), .C(N1257), .D(N1258), .Y(N218) );
  NAND4X1TF U1165 ( .A(N1259), .B(N1260), .C(N1261), .D(N1262), .Y(N217) );
  NAND4X1TF U1166 ( .A(N1263), .B(N1264), .C(N1265), .D(N1266), .Y(N216) );
  NAND4X1TF U1167 ( .A(N1267), .B(N1268), .C(N1269), .D(N1270), .Y(N215) );
  NAND4X1TF U1168 ( .A(N1271), .B(N1272), .C(N1273), .D(N1274), .Y(N214) );
  NAND4X1TF U1169 ( .A(N1275), .B(N1276), .C(N1277), .D(N1278), .Y(N213) );
  NAND4X1TF U1170 ( .A(N1279), .B(N1280), .C(N1281), .D(N1282), .Y(N212) );
  NAND4X1TF U1171 ( .A(N1283), .B(N1284), .C(N1285), .D(N1286), .Y(N211) );
  NAND4X1TF U1172 ( .A(N1287), .B(N1288), .C(N1289), .D(N1290), .Y(N210) );
  NAND4X1TF U1173 ( .A(N1291), .B(N1292), .C(N1293), .D(N1294), .Y(N209) );
  NAND4X1TF U1174 ( .A(N1295), .B(N1296), .C(N1297), .D(N1298), .Y(N208) );
  NAND4X1TF U1175 ( .A(N1299), .B(N1300), .C(N1301), .D(N1302), .Y(N207) );
  NAND4X1TF U1176 ( .A(N1311), .B(N1312), .C(N1313), .D(N1314), .Y(N262) );
  NAND4X1TF U1177 ( .A(N1315), .B(N1316), .C(N1317), .D(N1318), .Y(N261) );
  NAND4X1TF U1178 ( .A(N1319), .B(N1320), .C(N1321), .D(N1322), .Y(N260) );
  NAND4X1TF U1179 ( .A(N1323), .B(N1324), .C(N1325), .D(N1326), .Y(N259) );
  NAND4X1TF U1180 ( .A(N1327), .B(N1328), .C(N1329), .D(N1330), .Y(N258) );
  NAND4X1TF U1181 ( .A(N1331), .B(N1332), .C(N1333), .D(N1334), .Y(N257) );
  NAND4X1TF U1182 ( .A(N1335), .B(N1336), .C(N1337), .D(N1338), .Y(N256) );
  NAND4X1TF U1183 ( .A(N1339), .B(N1340), .C(N1341), .D(N1342), .Y(N255) );
  NAND4X1TF U1184 ( .A(N1343), .B(N1344), .C(N1345), .D(N1346), .Y(N254) );
  NAND4X1TF U1185 ( .A(N1347), .B(N1348), .C(N1349), .D(N1350), .Y(N253) );
  NAND4X1TF U1186 ( .A(N1351), .B(N1352), .C(N1353), .D(N1354), .Y(N252) );
  NAND4X1TF U1187 ( .A(N1355), .B(N1356), .C(N1357), .D(N1358), .Y(N251) );
  NAND4X1TF U1188 ( .A(N1359), .B(N1360), .C(N1361), .D(N1362), .Y(N250) );
  NAND4X1TF U1189 ( .A(N1363), .B(N1364), .C(N1365), .D(N1366), .Y(N249) );
  NAND4X1TF U1190 ( .A(N1367), .B(N1368), .C(N1369), .D(N1370), .Y(N248) );
  NAND4X1TF U1191 ( .A(N1371), .B(N1372), .C(N1373), .D(N1374), .Y(N247) );
endmodule


module SCPU_SRAM_8BIT_ALU_SPI_TOP_VG ( CLK, RST_N, CTRL_MODE, CTRL_BGN, CPU_BGN, 
        LOAD_N, CTRL_SI, APP_DONE, ADC_PI, TEST_MUX, CPU_WAIT, CTRL_RDY, 
        APP_START, CTRL_SO, NXT, SCLK1, SCLK2, LAT, SPI_SO );
  input [1:0] CTRL_MODE;
  input [9:0] ADC_PI;
  input [2:0] TEST_MUX;
  output [1:0] NXT;
  input CLK, RST_N, CTRL_BGN, CPU_BGN, LOAD_N, CTRL_SI, APP_DONE, CPU_WAIT;
  output CTRL_RDY, APP_START, CTRL_SO, SCLK1, SCLK2, LAT, SPI_SO;
  wire   CEN_AFTER_MUX, WEN_AFTER_MUX, I_CLK, I_RST_N, I_CTRL_BGN, I_CPU_BGN,
         I_LOAD_N, I_CTRL_SI, I_APP_DONE, I_CPU_WAIT, I_APP_START, I_CTRL_SO,
         I_SCLK1, I_SCLK2, I_LAT, I_SPI_SO, SCPU_CTRL_SPI_I_SPI_SO,
         \SCPU_CTRL_SPI_POUT[0] , \SCPU_CTRL_SPI_POUT[1] ,
         \SCPU_CTRL_SPI_POUT[2] , \SCPU_CTRL_SPI_POUT[3] ,
         \SCPU_CTRL_SPI_POUT[4] , \SCPU_CTRL_SPI_POUT[5] ,
         \SCPU_CTRL_SPI_POUT[6] , \SCPU_CTRL_SPI_POUT[7] ,
         \SCPU_CTRL_SPI_POUT[8] , \SCPU_CTRL_SPI_POUT[9] ,
         \SCPU_CTRL_SPI_POUT[10] , \SCPU_CTRL_SPI_POUT[11] ,
         \SCPU_CTRL_SPI_POUT[12] , \SCPU_CTRL_SPI_FOUT[0] ,
         \SCPU_CTRL_SPI_FOUT[1] , \SCPU_CTRL_SPI_FOUT[2] ,
         \SCPU_CTRL_SPI_FOUT[3] , \SCPU_CTRL_SPI_FOUT[4] ,
         \SCPU_CTRL_SPI_FOUT[5] , \SCPU_CTRL_SPI_FOUT[6] ,
         \SCPU_CTRL_SPI_FOUT[7] , \SCPU_CTRL_SPI_FOUT[8] ,
         \SCPU_CTRL_SPI_FOUT[9] , \SCPU_CTRL_SPI_FOUT[10] ,
         \SCPU_CTRL_SPI_FOUT[11] , \SCPU_CTRL_SPI_FOUT[12] , SCPU_CTRL_SPI_CEN,
         \SCPU_CTRL_SPI_IO_DATAOUTB[0] , \SCPU_CTRL_SPI_IO_DATAOUTB[1] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[2] , \SCPU_CTRL_SPI_IO_DATAOUTB[3] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[4] , \SCPU_CTRL_SPI_IO_DATAOUTB[5] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[6] , \SCPU_CTRL_SPI_IO_DATAOUTB[7] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[8] , \SCPU_CTRL_SPI_IO_DATAOUTB[9] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[10] , \SCPU_CTRL_SPI_IO_DATAOUTB[11] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[12] , \SCPU_CTRL_SPI_IO_DATAOUTA[0] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[1] , \SCPU_CTRL_SPI_IO_DATAOUTA[2] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[3] , \SCPU_CTRL_SPI_IO_DATAOUTA[4] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[5] , \SCPU_CTRL_SPI_IO_DATAOUTA[6] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[7] , \SCPU_CTRL_SPI_IO_DATAOUTA[8] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[9] , \SCPU_CTRL_SPI_IO_DATAOUTA[10] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[11] , \SCPU_CTRL_SPI_IO_DATAOUTA[12] ,
         \SCPU_CTRL_SPI_IO_DATAINA[0] , \SCPU_CTRL_SPI_IO_DATAINA[1] ,
         \SCPU_CTRL_SPI_IO_DATAINA[2] , \SCPU_CTRL_SPI_IO_DATAINA[3] ,
         \SCPU_CTRL_SPI_IO_DATAINA[4] , \SCPU_CTRL_SPI_IO_DATAINA[5] ,
         \SCPU_CTRL_SPI_IO_DATAINA[6] , \SCPU_CTRL_SPI_IO_DATAINA[7] ,
         \SCPU_CTRL_SPI_IO_DATAINA[8] , \SCPU_CTRL_SPI_IO_DATAINA[9] ,
         \SCPU_CTRL_SPI_IO_DATAINA[10] , \SCPU_CTRL_SPI_IO_DATAINA[11] ,
         \SCPU_CTRL_SPI_IO_DATAINA[12] , SCPU_CTRL_SPI_IO_CONTROL_0,
         SCPU_CTRL_SPI_IO_CONTROL_1, SCPU_CTRL_SPI_IO_CONTROL_2,
         SCPU_CTRL_SPI_IO_CONTROL_3, SCPU_CTRL_SPI_IO_CONTROL_4,
         SCPU_CTRL_SPI_IO_CONTROL_5, SCPU_CTRL_SPI_IO_CONTROL_6,
         \SCPU_CTRL_SPI_IO_STATUS[0] , SCPU_CTRL_SPI_D_WE,
         SCPU_CTRL_SPI_IS_I_ADDR, SCPU_CTRL_SPI_CCT_N57, SCPU_CTRL_SPI_CCT_N56,
         SCPU_CTRL_SPI_CCT_N55, SCPU_CTRL_SPI_CCT_N53, SCPU_CTRL_SPI_CCT_N52,
         SCPU_CTRL_SPI_CCT_IS_SHIFT, \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[3] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[5] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[7] , \SCPU_CTRL_SPI_CCT_REG_BITS[1] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[2] , \SCPU_CTRL_SPI_CCT_REG_BITS[3] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[4] , \SCPU_CTRL_SPI_CCT_REG_BITS[5] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[6] , \SCPU_CTRL_SPI_CCT_REG_BITS[7] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[8] , \SCPU_CTRL_SPI_CCT_REG_BITS[9] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[10] , \SCPU_CTRL_SPI_CCT_REG_BITS[11] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[12] , \SCPU_CTRL_SPI_CCT_REG_BITS[13] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[14] , \SCPU_CTRL_SPI_CCT_REG_BITS[15] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[16] , \SCPU_CTRL_SPI_CCT_REG_BITS[17] ,
         \SCPU_CTRL_SPI_CCT_CTRL_STATE[0] , SCPU_CTRL_SPI_PUT_N112,
         SCPU_CTRL_SPI_PUT_N111, SCPU_CTRL_SPI_PUT_N110,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] , SCPU_CTRL_SPI_PUT_N27,
         SCPU_CTRL_SPI_PUT_IS_ADDR_LEN_NZ, \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ,
         \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ,
         \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] ,
         \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[4] , \SCPU_CTRL_SPI_PUT_SPI_STATE[1] ,
         \SCPU_CTRL_SPI_PUT_CNT_STATE[0] , \SCPU_CTRL_SPI_PUT_CNT_STATE[1] ,
         \SCPU_CTRL_SPI_PUT_CNT_STATE[2] , N34, N35, N36, N37, N38, N39, N40,
         N41, N42, N43, N44, N45, N46, N47, N48, N87, N88, N89, N90, N91, N92,
         N93, N94, N95, N96, N100, N102, N108, N110, N111, N168, N174, N175,
         N233, N234, N235, N236, N237, N238, N239, N240, N241, N242, N243,
         N244, N245, N246, N247, N248, N249, N250, N251, N252, N253, N254,
         N256, N257, N258, N259, N260, N261, N263, N264, N265, N266, N277,
         N278, N279, N280, N281, N282, N283, N311, N312, N313, N314, N315,
         N316, N317, N318, N319, N320, N323, N324, N325, N326, N327, N328,
         N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, N339,
         N340, N341, N342, N343, N344, N345, N346, N347, N348, N349, N350,
         N351, N352, N353, N354, N355, N356, N357, N358, N359, N360, N361,
         N362, N363, N364, N365, N366, N367, N368, N369, N370, N371, N372,
         N373, N374, N375, N376, N377, N378, N379, N380, N381, N382, N383,
         N384, N385, N386, N387, N388, N389, N390, N391, N392, N393, N394,
         N395, N396, N397, N398, N399, N400, N401, N402, N403, N404, N405,
         N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416,
         N417, N418, N419, N420, N421, N422, N423, N424, N425, N426, N427,
         N428, N429, N430, N431, N432, N433, N434, N435, N436, N437, N438,
         N439, N440, N441, N442, N443, N444, N445, N446, N447, N448, N449,
         N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460,
         N461, N462, N463, N464, N465, N466, N467, N468, N469, N470, N471,
         N472, N473, N474, N475, N476, N477, N478, N479, N480, N481, N482,
         N483, N484, N485, N486, N487, N488, N489, N490, N491, N492, N493,
         N494, N495, N496, N497, N498, N499, N500, N501, N502, N503, N504,
         N505, N506, N507, N508, N509, N510, N511, N512, N513, N514, N515,
         N516;
  wire   [9:0] A_AFTER_MUX;
  wire   [7:0] D_AFTER_MUX;
  wire   [7:0] Q_FROM_SRAM;
  wire   [1:0] I_CTRL_MODE;
  wire   [9:0] I_ADC_PI;
  wire   [2:0] I_TEST_MUX;
  wire   [1:0] I_NXT;
  wire   [9:0] SCPU_CTRL_SPI_A_SPI;
  wire   [9:0] SCPU_CTRL_SPI_IO_OFFSET;
  wire   [7:0] SCPU_CTRL_SPI_D_DATAOUT;
  wire   [9:1] SCPU_CTRL_SPI_D_ADDR;
  wire   [9:0] SCPU_CTRL_SPI_I_ADDR;
  wire   [1:0] SCPU_CTRL_SPI_I_NXT;
  wire   [7:0] SCPU_CTRL_SPI_D_DATAIN;
  wire   [7:0] SCPU_CTRL_SPI_I_DATAIN;
  wire   [7:1] SCPU_CTRL_SPI_PUT_SRAM_REGS;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12;

  RA1SHD_IBM1024X8 sram ( .Q(Q_FROM_SRAM), .A(A_AFTER_MUX), .D(D_AFTER_MUX), 
        .CLK(I_CLK), .CEN(CEN_AFTER_MUX), .WEN(WEN_AFTER_MUX) );
  PIC ipad_clk ( .IE(1'b1), .P(CLK), .Y(I_CLK) );
  PIC ipad_rst_n ( .IE(1'b1), .P(RST_N), .Y(I_RST_N) );
  PIC ipad_ctrl_mode0 ( .IE(1'b1), .P(CTRL_MODE[0]), .Y(I_CTRL_MODE[0]) );
  PIC ipad_ctrl_mode1 ( .IE(1'b1), .P(CTRL_MODE[1]), .Y(I_CTRL_MODE[1]) );
  PIC ipad_ctrl_bgn ( .IE(1'b1), .P(CTRL_BGN), .Y(I_CTRL_BGN) );
  PIC ipad_cpu_bgn ( .IE(1'b1), .P(CPU_BGN), .Y(I_CPU_BGN) );
  PIC ipad_load_n ( .IE(1'b1), .P(LOAD_N), .Y(I_LOAD_N) );
  PIC ipad_ctrl_si ( .IE(1'b1), .P(CTRL_SI), .Y(I_CTRL_SI) );
  PIC ipad_app_done ( .IE(1'b1), .P(APP_DONE), .Y(I_APP_DONE) );
  PIC ipad_adc_pi0 ( .IE(1'b1), .P(ADC_PI[0]), .Y(I_ADC_PI[0]) );
  PIC ipad_adc_pi1 ( .IE(1'b1), .P(ADC_PI[1]), .Y(I_ADC_PI[1]) );
  PIC ipad_adc_pi2 ( .IE(1'b1), .P(ADC_PI[2]), .Y(I_ADC_PI[2]) );
  PIC ipad_adc_pi3 ( .IE(1'b1), .P(ADC_PI[3]), .Y(I_ADC_PI[3]) );
  PIC ipad_adc_pi4 ( .IE(1'b1), .P(ADC_PI[4]), .Y(I_ADC_PI[4]) );
  PIC ipad_adc_pi5 ( .IE(1'b1), .P(ADC_PI[5]), .Y(I_ADC_PI[5]) );
  PIC ipad_adc_pi6 ( .IE(1'b1), .P(ADC_PI[6]), .Y(I_ADC_PI[6]) );
  PIC ipad_adc_pi7 ( .IE(1'b1), .P(ADC_PI[7]), .Y(I_ADC_PI[7]) );
  PIC ipad_adc_pi8 ( .IE(1'b1), .P(ADC_PI[8]), .Y(I_ADC_PI[8]) );
  PIC ipad_adc_pi9 ( .IE(1'b1), .P(ADC_PI[9]), .Y(I_ADC_PI[9]) );
  PIC ipad_test_mux0 ( .IE(1'b1), .P(TEST_MUX[0]), .Y(I_TEST_MUX[0]) );
  PIC ipad_test_mux1 ( .IE(1'b1), .P(TEST_MUX[1]), .Y(I_TEST_MUX[1]) );
  PIC ipad_test_mux2 ( .IE(1'b1), .P(TEST_MUX[2]), .Y(I_TEST_MUX[2]) );
  PIC ipad_cpu_wait ( .IE(1'b1), .P(CPU_WAIT), .Y(I_CPU_WAIT) );
  POC8B opad_app_start ( .A(I_APP_START), .P(APP_START) );
  POC8B opad_ctrl_rdy ( .A(N265), .P(CTRL_RDY) );
  POC8B opad_ctrl_so ( .A(I_CTRL_SO), .P(CTRL_SO) );
  POC8B opad_nxt0 ( .A(I_NXT[0]), .P(NXT[0]) );
  POC8B opad_nxt1 ( .A(I_NXT[1]), .P(NXT[1]) );
  POC8B opad_sclk1 ( .A(I_SCLK1), .P(SCLK1) );
  POC8B opad_sclk2 ( .A(I_SCLK2), .P(SCLK2) );
  POC8B opad_lat ( .A(I_LAT), .P(LAT) );
  POC8B opad_spi_so ( .A(I_SPI_SO), .P(SPI_SO) );
  SHARE_SUPERALU_VG \scpu_ctrl_spi/ALU_01  ( .CLK(I_CLK), .RST_N(I_RST_N), .X_IN(
        {\SCPU_CTRL_SPI_IO_DATAOUTA[12] , \SCPU_CTRL_SPI_IO_DATAOUTA[11] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[10] , \SCPU_CTRL_SPI_IO_DATAOUTA[9] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[8] , \SCPU_CTRL_SPI_IO_DATAOUTA[7] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[6] , \SCPU_CTRL_SPI_IO_DATAOUTA[5] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[4] , \SCPU_CTRL_SPI_IO_DATAOUTA[3] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[2] , \SCPU_CTRL_SPI_IO_DATAOUTA[1] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[0] }), .Y_IN({
        \SCPU_CTRL_SPI_IO_DATAOUTB[12] , \SCPU_CTRL_SPI_IO_DATAOUTB[11] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[10] , \SCPU_CTRL_SPI_IO_DATAOUTB[9] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[8] , \SCPU_CTRL_SPI_IO_DATAOUTB[7] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[6] , \SCPU_CTRL_SPI_IO_DATAOUTB[5] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[4] , \SCPU_CTRL_SPI_IO_DATAOUTB[3] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[2] , \SCPU_CTRL_SPI_IO_DATAOUTB[1] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[0] }), .ALU_START(N318), .ALU_TYPE({
        SCPU_CTRL_SPI_IO_CONTROL_4, SCPU_CTRL_SPI_IO_CONTROL_3, 
        SCPU_CTRL_SPI_IO_CONTROL_2}), .MODE_TYPE({SCPU_CTRL_SPI_IO_CONTROL_1, 
        SCPU_CTRL_SPI_IO_CONTROL_0}), .OFFSET(SCPU_CTRL_SPI_IO_OFFSET), .FOUT(
        {\SCPU_CTRL_SPI_FOUT[12] , \SCPU_CTRL_SPI_FOUT[11] , 
        \SCPU_CTRL_SPI_FOUT[10] , \SCPU_CTRL_SPI_FOUT[9] , 
        \SCPU_CTRL_SPI_FOUT[8] , \SCPU_CTRL_SPI_FOUT[7] , 
        \SCPU_CTRL_SPI_FOUT[6] , \SCPU_CTRL_SPI_FOUT[5] , 
        \SCPU_CTRL_SPI_FOUT[4] , \SCPU_CTRL_SPI_FOUT[3] , 
        \SCPU_CTRL_SPI_FOUT[2] , \SCPU_CTRL_SPI_FOUT[1] , 
        \SCPU_CTRL_SPI_FOUT[0] }), .POUT({\SCPU_CTRL_SPI_POUT[12] , 
        \SCPU_CTRL_SPI_POUT[11] , \SCPU_CTRL_SPI_POUT[10] , 
        \SCPU_CTRL_SPI_POUT[9] , \SCPU_CTRL_SPI_POUT[8] , 
        \SCPU_CTRL_SPI_POUT[7] , \SCPU_CTRL_SPI_POUT[6] , 
        \SCPU_CTRL_SPI_POUT[5] , \SCPU_CTRL_SPI_POUT[4] , 
        \SCPU_CTRL_SPI_POUT[3] , \SCPU_CTRL_SPI_POUT[2] , 
        \SCPU_CTRL_SPI_POUT[1] , \SCPU_CTRL_SPI_POUT[0] }), .ALU_IS_DONE(
        \SCPU_CTRL_SPI_IO_STATUS[0] ) );
  SERIAL_CPU_8BIT_VG \scpu_ctrl_spi/uut  ( .CLK(I_CLK), .ENABLE(1'b0), .RST_N(
        I_RST_N), .START(I_CPU_BGN), .I_DATAIN(SCPU_CTRL_SPI_I_DATAIN), 
        .D_DATAIN(SCPU_CTRL_SPI_D_DATAIN), .CPU_WAIT(I_CPU_WAIT), .IS_I_ADDR(
        SCPU_CTRL_SPI_IS_I_ADDR), .NXT(SCPU_CTRL_SPI_I_NXT), .I_ADDR(
        SCPU_CTRL_SPI_I_ADDR), .D_ADDR({SCPU_CTRL_SPI_D_ADDR, 
        SYNOPSYS_UNCONNECTED__0}), .D_WE(SCPU_CTRL_SPI_D_WE), .D_DATAOUT(
        SCPU_CTRL_SPI_D_DATAOUT), .IO_STATUS({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, I_APP_DONE, N266, 
        \SCPU_CTRL_SPI_IO_STATUS[0] }), .IO_DATAINA({1'b0, 1'b0, 1'b0, 
        \SCPU_CTRL_SPI_IO_DATAINA[12] , \SCPU_CTRL_SPI_IO_DATAINA[11] , 
        \SCPU_CTRL_SPI_IO_DATAINA[10] , \SCPU_CTRL_SPI_IO_DATAINA[9] , 
        \SCPU_CTRL_SPI_IO_DATAINA[8] , \SCPU_CTRL_SPI_IO_DATAINA[7] , 
        \SCPU_CTRL_SPI_IO_DATAINA[6] , \SCPU_CTRL_SPI_IO_DATAINA[5] , 
        \SCPU_CTRL_SPI_IO_DATAINA[4] , \SCPU_CTRL_SPI_IO_DATAINA[3] , 
        \SCPU_CTRL_SPI_IO_DATAINA[2] , \SCPU_CTRL_SPI_IO_DATAINA[1] , 
        \SCPU_CTRL_SPI_IO_DATAINA[0] }), .IO_DATAINB({1'b0, 1'b0, 1'b0, 
        \SCPU_CTRL_SPI_POUT[12] , \SCPU_CTRL_SPI_POUT[11] , 
        \SCPU_CTRL_SPI_POUT[10] , \SCPU_CTRL_SPI_POUT[9] , 
        \SCPU_CTRL_SPI_POUT[8] , \SCPU_CTRL_SPI_POUT[7] , 
        \SCPU_CTRL_SPI_POUT[6] , \SCPU_CTRL_SPI_POUT[5] , 
        \SCPU_CTRL_SPI_POUT[4] , \SCPU_CTRL_SPI_POUT[3] , 
        \SCPU_CTRL_SPI_POUT[2] , \SCPU_CTRL_SPI_POUT[1] , 
        \SCPU_CTRL_SPI_POUT[0] }), .IO_DATAOUTA({SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        \SCPU_CTRL_SPI_IO_DATAOUTA[12] , \SCPU_CTRL_SPI_IO_DATAOUTA[11] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[10] , \SCPU_CTRL_SPI_IO_DATAOUTA[9] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[8] , \SCPU_CTRL_SPI_IO_DATAOUTA[7] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[6] , \SCPU_CTRL_SPI_IO_DATAOUTA[5] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[4] , \SCPU_CTRL_SPI_IO_DATAOUTA[3] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[2] , \SCPU_CTRL_SPI_IO_DATAOUTA[1] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[0] }), .IO_DATAOUTB({
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, \SCPU_CTRL_SPI_IO_DATAOUTB[12] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[11] , \SCPU_CTRL_SPI_IO_DATAOUTB[10] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[9] , \SCPU_CTRL_SPI_IO_DATAOUTB[8] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[7] , \SCPU_CTRL_SPI_IO_DATAOUTB[6] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[5] , \SCPU_CTRL_SPI_IO_DATAOUTB[4] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[3] , \SCPU_CTRL_SPI_IO_DATAOUTB[2] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[1] , \SCPU_CTRL_SPI_IO_DATAOUTB[0] }), 
        .IO_OFFSET({SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SCPU_CTRL_SPI_IO_OFFSET}), .\IO_CONTROL[7] (I_APP_START), 
        .\IO_CONTROL[6] (SCPU_CTRL_SPI_IO_CONTROL_6), .\IO_CONTROL[5]_BAR (
        SCPU_CTRL_SPI_IO_CONTROL_5), .\IO_CONTROL[4] (
        SCPU_CTRL_SPI_IO_CONTROL_4), .\IO_CONTROL[3] (
        SCPU_CTRL_SPI_IO_CONTROL_3), .\IO_CONTROL[2] (
        SCPU_CTRL_SPI_IO_CONTROL_2), .\IO_CONTROL[1] (
        SCPU_CTRL_SPI_IO_CONTROL_1), .\IO_CONTROL[0] (
        SCPU_CTRL_SPI_IO_CONTROL_0) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[7]  ( .D(N168), .RN(
        SCPU_CTRL_SPI_CCT_N57), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[7] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[5]  ( .D(N168), .RN(
        SCPU_CTRL_SPI_CCT_N55), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[5] ), .QN(N335) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[3]  ( .D(N168), .RN(
        SCPU_CTRL_SPI_CCT_N53), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[3] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[2]  ( .D(N168), .RN(
        SCPU_CTRL_SPI_CCT_N52), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ), .QN(N337) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[6]  ( .D(N168), .RN(
        SCPU_CTRL_SPI_CCT_N56), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[17]  ( .D(I_CTRL_SI), .E(N344), 
        .CK(I_CLK), .Q(\SCPU_CTRL_SPI_CCT_REG_BITS[17] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[16]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[17] ), .E(N344), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[16] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[15]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[16] ), .E(N100), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[15] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[14]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[15] ), .E(N100), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[14] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[13]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[14] ), .E(N100), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[13] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[12]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[13] ), .E(N100), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[12] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[11]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[12] ), .E(N100), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[11] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[10]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[11] ), .E(N100), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[10] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[9]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[10] ), .E(N100), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[9] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[8]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[9] ), .E(N100), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[8] ) );
  DFFSX2TF \scpu_ctrl_spi/put/cnt_state_reg[0]  ( .D(SCPU_CTRL_SPI_PUT_N110), 
        .CK(I_CLK), .SN(SCPU_CTRL_SPI_IO_CONTROL_6), .Q(
        \SCPU_CTRL_SPI_PUT_CNT_STATE[0] ), .QN(N336) );
  DFFRX2TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[3]  ( .D(N252), .CK(I_CLK), 
        .RN(N317), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ), .QN(N340) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[2]  ( .D(N42), .CK(I_CLK), 
        .SN(N41), .RN(N40), .QN(N339) );
  DFFRX2TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[0]  ( .D(N249), .CK(I_CLK), 
        .RN(N317), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .QN(N334) );
  DFFRX2TF \scpu_ctrl_spi/put/spi_state_reg[0]  ( .D(N253), .CK(I_CLK), .RN(
        N317), .Q(N330), .QN(N108) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[4]  ( .D(N48), .CK(I_CLK), 
        .SN(N47), .RN(N46), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[4] ), .QN(N328)
         );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[1]  ( .D(N39), .CK(I_CLK), 
        .SN(N38), .RN(N37), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ), .QN(N326)
         );
  DFFRX2TF \scpu_ctrl_spi/put/cnt_state_reg[1]  ( .D(SCPU_CTRL_SPI_PUT_N111), 
        .CK(I_CLK), .RN(N317), .Q(\SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .QN(N325)
         );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[3]  ( .D(N45), .CK(I_CLK), 
        .SN(N44), .RN(N43), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] ), .QN(N324)
         );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[7]  ( .D(N248), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[7]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[6]  ( .D(N242), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[6]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[5]  ( .D(N243), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[5]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[4]  ( .D(N244), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[4]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[3]  ( .D(N245), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[3]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[2]  ( .D(N246), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[2]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[1]  ( .D(N247), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[1]) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[7]  ( .D(N233), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[7] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[6]  ( .D(N234), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[6] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[5]  ( .D(N235), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[5] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[4]  ( .D(N236), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[4] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[3]  ( .D(N237), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[3] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[2]  ( .D(N238), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[2] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[1]  ( .D(N239), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[1] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/is_shift_reg  ( .D(N174), .RN(N175), .CK(I_CLK), 
        .QN(SCPU_CTRL_SPI_CCT_IS_SHIFT) );
  DFFQX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[1]  ( .D(N258), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[4]  ( .D(N260), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[0]  ( .D(N259), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[0]  ( .D(N240), .CK(I_CLK), .Q(
        I_CTRL_SO) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[0]  ( .D(N241), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_I_SPI_SO) );
  DFFXLTF \scpu_ctrl_spi/cct/ctrl_state_reg[0]  ( .D(N261), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .QN(N341) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[0]  ( .D(N36), .CK(I_CLK), 
        .SN(N35), .RN(N34), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ) );
  DFFRX2TF \scpu_ctrl_spi/put/spi_state_reg[2]  ( .D(N256), .CK(I_CLK), .RN(
        N317), .Q(N323), .QN(N110) );
  DFFNSRX4TF \scpu_ctrl_spi/put/spi_MUX_reg  ( .D(N257), .CKN(I_CLK), .SN(1'b1), .RN(1'b1), .Q(N342), .QN(N111) );
  DFFNSRXLTF \scpu_ctrl_spi/cct/CEN_reg  ( .D(N264), .CKN(I_CLK), .SN(1'b1), 
        .RN(1'b1), .Q(SCPU_CTRL_SPI_CEN) );
  DFFNSRXLTF \scpu_ctrl_spi/put/is_addr_len_nz_reg  ( .D(SCPU_CTRL_SPI_PUT_N27), .CKN(I_CLK), .SN(1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_PUT_IS_ADDR_LEN_NZ) );
  DFFNSRXLTF \scpu_ctrl_spi/put/sram_addr_reg[9]  ( .D(N96), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[9]) );
  EDFFTRXLTF \scpu_ctrl_spi/cct/ctrl_state_reg[1]  ( .RN(I_CTRL_BGN), .D(1'b1), 
        .E(N283), .CK(I_CLK), .Q(N327), .QN(N102) );
  DFFRX1TF \scpu_ctrl_spi/put/cnt_state_reg[2]  ( .D(SCPU_CTRL_SPI_PUT_N112), 
        .CK(I_CLK), .RN(N317), .Q(\SCPU_CTRL_SPI_PUT_CNT_STATE[2] ) );
  DFFRX1TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[1]  ( .D(N250), .CK(I_CLK), 
        .RN(N317), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ) );
  DFFRX1TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[2]  ( .D(N251), .CK(I_CLK), 
        .RN(N316), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ) );
  DFFRX2TF \scpu_ctrl_spi/put/spi_state_reg[1]  ( .D(N254), .CK(I_CLK), .RN(
        N317), .Q(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[1]  ( .D(N88), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[1]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[3]  ( .D(N90), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[3]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[2]  ( .D(N89), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[2]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[6]  ( .D(N93), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[6]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[4]  ( .D(N91), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[4]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[7]  ( .D(N94), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[7]), .QN(N331) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[8]  ( .D(N95), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[8]), .QN(N333) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[0]  ( .D(N87), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[0]), .QN(N332) );
  DFFNSRX2TF \scpu_ctrl_spi/cct/D_WE_reg  ( .D(N263), .CKN(I_CLK), .SN(1'b1), 
        .RN(1'b1), .QN(N329) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[5]  ( .D(N92), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[5]), .QN(N338) );
  NOR3BX2TF U290 ( .AN(N339), .B(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .C(
        \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ), .Y(N515) );
  INVX2TF U291 ( .A(SCPU_CTRL_SPI_IO_CONTROL_5), .Y(N311) );
  AND2X2TF U292 ( .A(N312), .B(N329), .Y(N370) );
  AOI22XLTF U293 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[16] ), .A1(N312), .B0(
        SCPU_CTRL_SPI_D_ADDR[8]), .B1(N368), .Y(N277) );
  AOI22X1TF U294 ( .A0(N366), .A1(SCPU_CTRL_SPI_I_ADDR[8]), .B0(N367), .B1(
        SCPU_CTRL_SPI_A_SPI[8]), .Y(N278) );
  NAND2X1TF U295 ( .A(N277), .B(N278), .Y(A_AFTER_MUX[8]) );
  AOI22X1TF U296 ( .A0(SCPU_CTRL_SPI_A_SPI[9]), .A1(N367), .B0(
        SCPU_CTRL_SPI_I_ADDR[9]), .B1(N366), .Y(N279) );
  AOI22XLTF U297 ( .A0(SCPU_CTRL_SPI_D_ADDR[9]), .A1(N368), .B0(N312), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[17] ), .Y(N280) );
  NAND2X1TF U298 ( .A(N279), .B(N280), .Y(A_AFTER_MUX[9]) );
  OAI22X1TF U299 ( .A0(SCPU_CTRL_SPI_PUT_IS_ADDR_LEN_NZ), .A1(N511), .B0(N423), 
        .B1(N323), .Y(N281) );
  AOI21X1TF U300 ( .A0(N423), .A1(N323), .B0(N281), .Y(N282) );
  AOI22X1TF U301 ( .A0(N425), .A1(N282), .B0(N110), .B1(N428), .Y(N256) );
  OA21XLTF U302 ( .A0(N319), .A1(I_CTRL_MODE[0]), .B0(N410), .Y(N283) );
  AOI22XLTF U303 ( .A0(SCPU_CTRL_SPI_A_SPI[3]), .A1(N367), .B0(
        SCPU_CTRL_SPI_I_ADDR[3]), .B1(N366), .Y(N357) );
  AOI22XLTF U304 ( .A0(SCPU_CTRL_SPI_A_SPI[1]), .A1(N367), .B0(
        SCPU_CTRL_SPI_I_ADDR[1]), .B1(N366), .Y(N353) );
  OR2X2TF U320 ( .A(SCPU_CTRL_SPI_CEN), .B(N439), .Y(N369) );
  INVX2TF U321 ( .A(I_TEST_MUX[1]), .Y(N374) );
  NAND2XLTF U322 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[4] ), .B(N347), .Y(N47) );
  NAND2XLTF U323 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[3] ), .B(N347), .Y(N44) );
  NAND2BXLTF U324 ( .AN(\SCPU_CTRL_SPI_IO_DATAOUTB[3] ), .B(N343), .Y(N43) );
  NAND2XLTF U325 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[2] ), .B(N347), .Y(N41) );
  NAND2BXLTF U326 ( .AN(\SCPU_CTRL_SPI_IO_DATAOUTB[2] ), .B(N343), .Y(N40) );
  NAND2XLTF U327 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[1] ), .B(N347), .Y(N38) );
  NAND2BXLTF U328 ( .AN(\SCPU_CTRL_SPI_IO_DATAOUTB[1] ), .B(N343), .Y(N37) );
  NAND2XLTF U329 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[0] ), .B(N347), .Y(N35) );
  NAND2BXLTF U330 ( .AN(\SCPU_CTRL_SPI_IO_DATAOUTB[0] ), .B(N347), .Y(N34) );
  NAND2BXLTF U331 ( .AN(\SCPU_CTRL_SPI_IO_DATAOUTB[4] ), .B(N343), .Y(N46) );
  AND3X2TF U332 ( .A(N316), .B(N516), .C(SCPU_CTRL_SPI_PUT_IS_ADDR_LEN_NZ), 
        .Y(N507) );
  OAI211XLTF U333 ( .A0(N427), .A1(N330), .B0(N323), .C0(N425), .Y(N426) );
  INVX2TF U334 ( .A(N343), .Y(N316) );
  CLKBUFX2TF U335 ( .A(\SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .Y(N319) );
  AOI32X1TF U336 ( .A0(N111), .A1(N439), .A2(SCPU_CTRL_SPI_D_WE), .B0(
        I_CTRL_BGN), .B1(N329), .Y(WEN_AFTER_MUX) );
  NAND2XLTF U337 ( .A(SCPU_CTRL_SPI_A_SPI[0]), .B(SCPU_CTRL_SPI_A_SPI[1]), .Y(
        N504) );
  INVX2TF U338 ( .A(SCPU_CTRL_SPI_IO_CONTROL_6), .Y(N343) );
  INVX2TF U339 ( .A(N369), .Y(N312) );
  INVX2TF U340 ( .A(N369), .Y(N313) );
  INVX2TF U341 ( .A(N507), .Y(N314) );
  INVX2TF U342 ( .A(N507), .Y(N315) );
  INVX2TF U343 ( .A(N343), .Y(N317) );
  INVX2TF U344 ( .A(SCPU_CTRL_SPI_IO_CONTROL_5), .Y(N318) );
  OAI211X1TF U345 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] ), .A1(
        \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[4] ), .B0(N516), .C0(N515), .Y(N514)
         );
  NAND4BX2TF U346 ( .AN(N264), .B(I_CTRL_BGN), .C(SCPU_CTRL_SPI_CCT_IS_SHIFT), 
        .D(N453), .Y(N463) );
  AOI32XLTF U347 ( .A0(N516), .A1(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] ), .A2(
        N515), .B0(N514), .B1(N324), .Y(N45) );
  NOR3X4TF U348 ( .A(N108), .B(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .C(N323), 
        .Y(N516) );
  INVX2TF U349 ( .A(I_CTRL_BGN), .Y(N320) );
  NOR3X4TF U350 ( .A(N441), .B(N440), .C(N346), .Y(N450) );
  INVX2TF U351 ( .A(I_CTRL_BGN), .Y(N439) );
  NOR3X2TF U352 ( .A(I_TEST_MUX[0]), .B(N374), .C(N372), .Y(N402) );
  NOR2X2TF U353 ( .A(I_TEST_MUX[1]), .B(N371), .Y(N403) );
  NOR2X1TF U354 ( .A(N427), .B(N442), .Y(N438) );
  NOR3XLTF U355 ( .A(N319), .B(N327), .C(N439), .Y(N414) );
  NAND2X1TF U356 ( .A(I_CTRL_BGN), .B(N413), .Y(N420) );
  NOR2X1TF U357 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[3] ), .B(N348), .Y(N174)
         );
  CLKBUFX2TF U358 ( .A(N100), .Y(N344) );
  NAND2X1TF U359 ( .A(N363), .B(N362), .Y(A_AFTER_MUX[6]) );
  NAND2X1TF U360 ( .A(N361), .B(N360), .Y(A_AFTER_MUX[5]) );
  NAND2X1TF U361 ( .A(N359), .B(N358), .Y(A_AFTER_MUX[4]) );
  NAND2X1TF U362 ( .A(N357), .B(N356), .Y(A_AFTER_MUX[3]) );
  NAND2X1TF U363 ( .A(N355), .B(N354), .Y(A_AFTER_MUX[2]) );
  NAND2X1TF U364 ( .A(N353), .B(N352), .Y(A_AFTER_MUX[1]) );
  NAND2X1TF U365 ( .A(N365), .B(N364), .Y(A_AFTER_MUX[7]) );
  NOR2X2TF U366 ( .A(N342), .B(N464), .Y(N368) );
  NAND2BX2TF U367 ( .AN(SCPU_CTRL_SPI_IS_I_ADDR), .B(N439), .Y(N464) );
  CLKBUFX2TF U368 ( .A(N509), .Y(N345) );
  NAND4X1TF U369 ( .A(N397), .B(N396), .C(N395), .D(N394), .Y(I_SCLK2) );
  NAND4X1TF U370 ( .A(N379), .B(N378), .C(N377), .D(N376), .Y(I_LAT) );
  NAND4X1TF U371 ( .A(N387), .B(N386), .C(N385), .D(N384), .Y(I_NXT[1]) );
  NAND4X1TF U372 ( .A(N383), .B(N382), .C(N381), .D(N380), .Y(I_NXT[0]) );
  NAND4X1TF U373 ( .A(N392), .B(N391), .C(N390), .D(N389), .Y(I_SCLK1) );
  NAND4X1TF U374 ( .A(N409), .B(N408), .C(N407), .D(N406), .Y(I_SPI_SO) );
  INVX2TF U375 ( .A(I_TEST_MUX[0]), .Y(N373) );
  INVX2TF U376 ( .A(I_TEST_MUX[2]), .Y(N372) );
  AO21X1TF U377 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[3] ), .A1(N348), .B0(
        N174), .Y(SCPU_CTRL_SPI_CCT_N53) );
  OAI2BB2XLTF U378 ( .B0(N478), .B1(N477), .A0N(
        \SCPU_CTRL_SPI_PUT_CNT_STATE[2] ), .A1N(N476), .Y(
        SCPU_CTRL_SPI_PUT_N112) );
  NAND2X1TF U379 ( .A(N516), .B(N510), .Y(N512) );
  NOR2X1TF U380 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ), .B(N349), .Y(N350)
         );
  NAND2X1TF U381 ( .A(N335), .B(N411), .Y(N349) );
  NAND3X1TF U382 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .B(N110), .C(N330), 
        .Y(N437) );
  NOR2X1TF U383 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ), .B(N412), .Y(N411)
         );
  NAND2X1TF U384 ( .A(N174), .B(N175), .Y(N413) );
  OR3X1TF U385 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ), .B(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .C(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ), .Y(N348) );
  AND3X2TF U386 ( .A(SCPU_CTRL_SPI_CCT_IS_SHIFT), .B(N102), .C(N319), .Y(N100)
         );
  OAI2BB2XLTF U387 ( .B0(N428), .B1(N479), .A0N(
        \SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .A1N(N426), .Y(N254) );
  NOR2X1TF U388 ( .A(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ), .B(N424), .Y(N427)
         );
  OAI2BB1X1TF U389 ( .A0N(N313), .A1N(\SCPU_CTRL_SPI_CCT_REG_BITS[8] ), .B0(
        N351), .Y(A_AFTER_MUX[0]) );
  OAI221XLTF U390 ( .A0(N111), .A1(SCPU_CTRL_SPI_A_SPI[0]), .B0(N342), .B1(
        SCPU_CTRL_SPI_I_ADDR[0]), .C0(N439), .Y(N351) );
  AO22X1TF U391 ( .A0(N370), .A1(I_CTRL_SO), .B0(SCPU_CTRL_SPI_D_DATAOUT[0]), 
        .B1(N439), .Y(D_AFTER_MUX[0]) );
  NOR2X2TF U392 ( .A(N342), .B(N472), .Y(N366) );
  NAND2X2TF U393 ( .A(SCPU_CTRL_SPI_IS_I_ADDR), .B(N439), .Y(N472) );
  NOR2X2TF U394 ( .A(I_CTRL_BGN), .B(N111), .Y(N367) );
  NAND2X1TF U395 ( .A(N319), .B(N327), .Y(N264) );
  NOR2X1TF U396 ( .A(N466), .B(N464), .Y(SCPU_CTRL_SPI_D_DATAIN[1]) );
  NOR2X1TF U397 ( .A(N469), .B(N464), .Y(SCPU_CTRL_SPI_D_DATAIN[4]) );
  NOR2X1TF U398 ( .A(N473), .B(N464), .Y(SCPU_CTRL_SPI_D_DATAIN[7]) );
  NOR2X1TF U399 ( .A(N470), .B(N464), .Y(SCPU_CTRL_SPI_D_DATAIN[5]) );
  NOR2X1TF U400 ( .A(N467), .B(N464), .Y(SCPU_CTRL_SPI_D_DATAIN[2]) );
  NOR2X1TF U401 ( .A(N471), .B(N464), .Y(SCPU_CTRL_SPI_D_DATAIN[6]) );
  NOR2X1TF U402 ( .A(N468), .B(N464), .Y(SCPU_CTRL_SPI_D_DATAIN[3]) );
  CLKBUFX2TF U403 ( .A(N343), .Y(N347) );
  CLKBUFX2TF U404 ( .A(N343), .Y(N346) );
  NAND2X1TF U405 ( .A(N516), .B(SCPU_CTRL_SPI_PUT_IS_ADDR_LEN_NZ), .Y(N479) );
  OAI21X1TF U406 ( .A0(N418), .A1(N337), .B0(N348), .Y(SCPU_CTRL_SPI_CCT_N52)
         );
  NOR2X1TF U407 ( .A(\SCPU_CTRL_SPI_PUT_CNT_STATE[0] ), .B(N475), .Y(
        SCPU_CTRL_SPI_PUT_N110) );
  OAI211X1TF U408 ( .A0(N438), .A1(N334), .B0(N437), .C0(N436), .Y(N249) );
  AOI31X1TF U409 ( .A0(N516), .A1(N515), .A2(N324), .B0(N328), .Y(N48) );
  OAI211X1TF U410 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .A1(N436), .B0(
        N437), .C0(N435), .Y(N250) );
  OAI21X1TF U411 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .A1(N478), .B0(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .Y(N435) );
  OAI31X1TF U412 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .A1(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .A2(N478), .B0(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ), .Y(N434) );
  AOI22X1TF U413 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ), .A1(N432), .B0(
        N433), .B1(N340), .Y(N252) );
  AOI21X1TF U414 ( .A0(N440), .A1(N424), .B0(N478), .Y(N432) );
  NOR2X1TF U415 ( .A(N441), .B(N438), .Y(N478) );
  OAI21X1TF U416 ( .A0(N411), .A1(N335), .B0(N349), .Y(SCPU_CTRL_SPI_CCT_N55)
         );
  OAI32X1TF U417 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ), .A1(
        \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .A2(N512), .B0(N513), .B1(N326), 
        .Y(N39) );
  AOI32X1TF U418 ( .A0(N513), .A1(N514), .A2(N326), .B0(N339), .B1(N514), .Y(
        N42) );
  NOR2X1TF U419 ( .A(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .B(N511), .Y(N513)
         );
  OAI21X1TF U420 ( .A0(N452), .A1(N471), .B0(N448), .Y(N242) );
  AOI22X1TF U421 ( .A0(N450), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[6]), .B0(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[7]), .B1(N449), .Y(N448) );
  OAI21X1TF U422 ( .A0(N468), .A1(N452), .B0(N445), .Y(N245) );
  AOI22X1TF U423 ( .A0(N450), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[3]), .B0(N449), 
        .B1(SCPU_CTRL_SPI_PUT_SRAM_REGS[4]), .Y(N445) );
  OAI21X1TF U424 ( .A0(N470), .A1(N452), .B0(N447), .Y(N243) );
  AOI22X1TF U425 ( .A0(N450), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[5]), .B0(N449), 
        .B1(SCPU_CTRL_SPI_PUT_SRAM_REGS[6]), .Y(N447) );
  OAI21X1TF U426 ( .A0(N469), .A1(N452), .B0(N446), .Y(N244) );
  AOI22X1TF U427 ( .A0(N450), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[4]), .B0(N449), 
        .B1(SCPU_CTRL_SPI_PUT_SRAM_REGS[5]), .Y(N446) );
  OAI21X1TF U428 ( .A0(N467), .A1(N452), .B0(N444), .Y(N246) );
  AOI22X1TF U429 ( .A0(N450), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[2]), .B0(N449), 
        .B1(SCPU_CTRL_SPI_PUT_SRAM_REGS[3]), .Y(N444) );
  OAI21X1TF U430 ( .A0(N466), .A1(N452), .B0(N443), .Y(N247) );
  AOI22X1TF U431 ( .A0(N450), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[1]), .B0(N449), 
        .B1(SCPU_CTRL_SPI_PUT_SRAM_REGS[2]), .Y(N443) );
  OAI21X1TF U432 ( .A0(N465), .A1(N452), .B0(N451), .Y(N241) );
  AOI22X1TF U433 ( .A0(SCPU_CTRL_SPI_I_SPI_SO), .A1(N450), .B0(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[1]), .B1(N449), .Y(N451) );
  NOR2X2TF U434 ( .A(N346), .B(N442), .Y(N449) );
  INVX2TF U435 ( .A(N442), .Y(N440) );
  NAND3X2TF U436 ( .A(N439), .B(N317), .C(N441), .Y(N452) );
  INVX2TF U437 ( .A(N437), .Y(N441) );
  OAI22X1TF U438 ( .A0(I_CTRL_MODE[1]), .A1(N417), .B0(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .B1(N420), .Y(N259) );
  OAI21X1TF U439 ( .A0(N421), .A1(N420), .B0(N419), .Y(N258) );
  AOI21X1TF U440 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .A1(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ), .B0(N418), .Y(N421) );
  NOR2X1TF U441 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ), .B(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .Y(N418) );
  OAI21X1TF U442 ( .A0(N415), .A1(N420), .B0(N419), .Y(N260) );
  NOR3BX1TF U443 ( .AN(N414), .B(I_LOAD_N), .C(N413), .Y(N416) );
  AOI21X1TF U444 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ), .A1(N412), .B0(
        N411), .Y(N415) );
  INVX2TF U445 ( .A(N174), .Y(N412) );
  INVX2TF U446 ( .A(N420), .Y(N168) );
  NOR4X1TF U447 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[7] ), .B(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ), .C(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[5] ), .D(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ), .Y(N175) );
  OAI21X1TF U448 ( .A0(N470), .A1(N463), .B0(N459), .Y(N235) );
  AOI22X1TF U449 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[6] ), .A1(N344), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[5] ), .B1(N461), .Y(N459) );
  OAI21X1TF U450 ( .A0(N473), .A1(N463), .B0(N462), .Y(N233) );
  AOI22X1TF U451 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[8] ), .A1(N344), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[7] ), .B1(N461), .Y(N462) );
  OAI21X1TF U452 ( .A0(N468), .A1(N463), .B0(N457), .Y(N237) );
  AOI22X1TF U453 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[4] ), .A1(N344), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[3] ), .B1(N461), .Y(N457) );
  OAI21X1TF U454 ( .A0(N471), .A1(N463), .B0(N460), .Y(N234) );
  AOI22X1TF U455 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[7] ), .A1(N344), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[6] ), .B1(N461), .Y(N460) );
  OAI21X1TF U456 ( .A0(N466), .A1(N463), .B0(N455), .Y(N239) );
  AOI22X1TF U457 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[2] ), .A1(N344), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[1] ), .B1(N461), .Y(N455) );
  OAI21X1TF U458 ( .A0(N469), .A1(N463), .B0(N458), .Y(N236) );
  AOI22X1TF U459 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[5] ), .A1(N344), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[4] ), .B1(N461), .Y(N458) );
  OAI21X1TF U460 ( .A0(N467), .A1(N463), .B0(N456), .Y(N238) );
  AOI22X1TF U461 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[3] ), .A1(N344), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[2] ), .B1(N461), .Y(N456) );
  OAI21X1TF U462 ( .A0(N465), .A1(N463), .B0(N454), .Y(N240) );
  AOI22X1TF U463 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[1] ), .A1(N344), .B0(
        I_CTRL_SO), .B1(N461), .Y(N454) );
  OAI211X4TF U464 ( .A0(N102), .A1(N453), .B0(N319), .C0(
        SCPU_CTRL_SPI_CCT_IS_SHIFT), .Y(N461) );
  INVX2TF U465 ( .A(I_CTRL_MODE[1]), .Y(N453) );
  NOR2X1TF U466 ( .A(N102), .B(N319), .Y(N265) );
  AND2X2TF U467 ( .A(SCPU_CTRL_SPI_CEN), .B(I_CTRL_BGN), .Y(CEN_AFTER_MUX) );
  AOI32X1TF U468 ( .A0(N430), .A1(N429), .A2(N479), .B0(N428), .B1(N429), .Y(
        N253) );
  OAI21X1TF U469 ( .A0(N323), .A1(N477), .B0(N330), .Y(N429) );
  INVX2TF U470 ( .A(N475), .Y(N477) );
  INVX2TF U471 ( .A(N428), .Y(N425) );
  INVX2TF U472 ( .A(N431), .Y(N424) );
  NOR3X1TF U473 ( .A(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ), .B(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .C(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .Y(N431) );
  AOI21X1TF U474 ( .A0(N323), .A1(N423), .B0(N475), .Y(N428) );
  NOR3X1TF U475 ( .A(\SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .B(
        \SCPU_CTRL_SPI_PUT_CNT_STATE[0] ), .C(\SCPU_CTRL_SPI_PUT_CNT_STATE[2] ), .Y(N475) );
  NOR2X1TF U476 ( .A(N471), .B(N472), .Y(SCPU_CTRL_SPI_I_DATAIN[6]) );
  NOR2X1TF U477 ( .A(N466), .B(N472), .Y(SCPU_CTRL_SPI_I_DATAIN[1]) );
  NOR2X1TF U478 ( .A(N469), .B(N472), .Y(SCPU_CTRL_SPI_I_DATAIN[4]) );
  NOR2X1TF U479 ( .A(N465), .B(N472), .Y(SCPU_CTRL_SPI_I_DATAIN[0]) );
  NOR2X1TF U480 ( .A(N467), .B(N472), .Y(SCPU_CTRL_SPI_I_DATAIN[2]) );
  NOR2X1TF U481 ( .A(N470), .B(N472), .Y(SCPU_CTRL_SPI_I_DATAIN[5]) );
  NOR2X1TF U482 ( .A(N468), .B(N472), .Y(SCPU_CTRL_SPI_I_DATAIN[3]) );
  NOR2X1TF U483 ( .A(N473), .B(N472), .Y(SCPU_CTRL_SPI_I_DATAIN[7]) );
  AND2X2TF U484 ( .A(N510), .B(N317), .Y(SCPU_CTRL_SPI_PUT_N27) );
  AOI22X1TF U485 ( .A0(SCPU_CTRL_SPI_D_ADDR[6]), .A1(N368), .B0(N312), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[14] ), .Y(N362) );
  AOI22X1TF U486 ( .A0(SCPU_CTRL_SPI_A_SPI[6]), .A1(N367), .B0(
        SCPU_CTRL_SPI_I_ADDR[6]), .B1(N366), .Y(N363) );
  AOI22X1TF U487 ( .A0(SCPU_CTRL_SPI_D_ADDR[5]), .A1(N368), .B0(N313), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[13] ), .Y(N360) );
  AOI22X1TF U488 ( .A0(SCPU_CTRL_SPI_A_SPI[5]), .A1(N367), .B0(
        SCPU_CTRL_SPI_I_ADDR[5]), .B1(N366), .Y(N361) );
  AOI22X1TF U489 ( .A0(SCPU_CTRL_SPI_D_ADDR[4]), .A1(N368), .B0(N313), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[12] ), .Y(N358) );
  AOI22X1TF U490 ( .A0(SCPU_CTRL_SPI_A_SPI[4]), .A1(N367), .B0(
        SCPU_CTRL_SPI_I_ADDR[4]), .B1(N366), .Y(N359) );
  AOI22X1TF U491 ( .A0(SCPU_CTRL_SPI_D_ADDR[3]), .A1(N368), .B0(N313), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[11] ), .Y(N356) );
  AOI22X1TF U492 ( .A0(SCPU_CTRL_SPI_D_ADDR[2]), .A1(N368), .B0(N313), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[10] ), .Y(N354) );
  AOI22X1TF U493 ( .A0(SCPU_CTRL_SPI_A_SPI[2]), .A1(N367), .B0(
        SCPU_CTRL_SPI_I_ADDR[2]), .B1(N366), .Y(N355) );
  AOI22X1TF U494 ( .A0(SCPU_CTRL_SPI_D_ADDR[1]), .A1(N368), .B0(N313), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[9] ), .Y(N352) );
  AOI22X1TF U495 ( .A0(N368), .A1(SCPU_CTRL_SPI_D_ADDR[7]), .B0(N312), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[15] ), .Y(N364) );
  AOI22X1TF U496 ( .A0(SCPU_CTRL_SPI_A_SPI[7]), .A1(N367), .B0(N366), .B1(
        SCPU_CTRL_SPI_I_ADDR[7]), .Y(N365) );
  NOR2X1TF U497 ( .A(N465), .B(N464), .Y(SCPU_CTRL_SPI_D_DATAIN[0]) );
  OAI32X1TF U498 ( .A0(N346), .A1(N111), .A2(N422), .B0(N511), .B1(N346), .Y(
        N257) );
  INVX2TF U499 ( .A(N516), .Y(N511) );
  NOR2X1TF U500 ( .A(N108), .B(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .Y(N422) );
  OAI21X1TF U501 ( .A0(N345), .A1(N332), .B0(N508), .Y(N87) );
  AOI22X1TF U502 ( .A0(N507), .A1(N332), .B0(\SCPU_CTRL_SPI_IO_DATAOUTA[0] ), 
        .B1(N346), .Y(N508) );
  AOI22X1TF U503 ( .A0(N486), .A1(N331), .B0(\SCPU_CTRL_SPI_IO_DATAOUTA[7] ), 
        .B1(N347), .Y(N487) );
  OAI21X1TF U504 ( .A0(SCPU_CTRL_SPI_A_SPI[5]), .A1(N494), .B0(N493), .Y(N92)
         );
  AOI22X1TF U505 ( .A0(SCPU_CTRL_SPI_A_SPI[5]), .A1(N492), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[5] ), .B1(N347), .Y(N493) );
  OAI21X1TF U506 ( .A0(N491), .A1(N315), .B0(N345), .Y(N492) );
  OAI31X1TF U507 ( .A0(SCPU_CTRL_SPI_A_SPI[3]), .A1(N315), .A2(N501), .B0(N500), .Y(N90) );
  AOI22X1TF U508 ( .A0(SCPU_CTRL_SPI_A_SPI[3]), .A1(N499), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[3] ), .B1(N346), .Y(N500) );
  OAI21X1TF U509 ( .A0(N498), .A1(N314), .B0(N345), .Y(N499) );
  OAI31X1TF U510 ( .A0(SCPU_CTRL_SPI_A_SPI[1]), .A1(N315), .A2(N332), .B0(N506), .Y(N88) );
  AOI22X1TF U511 ( .A0(SCPU_CTRL_SPI_A_SPI[1]), .A1(N505), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[1] ), .B1(N346), .Y(N506) );
  OAI21X1TF U512 ( .A0(SCPU_CTRL_SPI_A_SPI[0]), .A1(N314), .B0(N345), .Y(N505)
         );
  OAI31X1TF U513 ( .A0(SCPU_CTRL_SPI_A_SPI[2]), .A1(N315), .A2(N504), .B0(N503), .Y(N89) );
  AOI22X1TF U514 ( .A0(SCPU_CTRL_SPI_A_SPI[2]), .A1(N502), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[2] ), .B1(N346), .Y(N503) );
  AOI32X1TF U515 ( .A0(SCPU_CTRL_SPI_A_SPI[0]), .A1(N345), .A2(
        SCPU_CTRL_SPI_A_SPI[1]), .B0(N315), .B1(N345), .Y(N502) );
  OAI31X1TF U516 ( .A0(SCPU_CTRL_SPI_A_SPI[4]), .A1(N315), .A2(N497), .B0(N496), .Y(N91) );
  AOI22X1TF U517 ( .A0(SCPU_CTRL_SPI_A_SPI[4]), .A1(N495), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[4] ), .B1(N347), .Y(N496) );
  AOI32X1TF U518 ( .A0(N498), .A1(N345), .A2(SCPU_CTRL_SPI_A_SPI[3]), .B0(N315), .B1(N345), .Y(N495) );
  OAI31X1TF U519 ( .A0(SCPU_CTRL_SPI_A_SPI[6]), .A1(N338), .A2(N494), .B0(N490), .Y(N93) );
  AOI22X1TF U520 ( .A0(SCPU_CTRL_SPI_A_SPI[6]), .A1(N489), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[6] ), .B1(N347), .Y(N490) );
  AOI32X1TF U521 ( .A0(N491), .A1(N345), .A2(SCPU_CTRL_SPI_A_SPI[5]), .B0(N315), .B1(N345), .Y(N489) );
  OAI21X1TF U522 ( .A0(N485), .A1(N333), .B0(N484), .Y(N95) );
  OAI31X1TF U523 ( .A0(SCPU_CTRL_SPI_A_SPI[9]), .A1(N333), .A2(N483), .B0(N482), .Y(N96) );
  AOI22X1TF U524 ( .A0(SCPU_CTRL_SPI_A_SPI[9]), .A1(N481), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[9] ), .B1(N346), .Y(N482) );
  OAI21X1TF U525 ( .A0(SCPU_CTRL_SPI_A_SPI[8]), .A1(N315), .B0(N485), .Y(N481)
         );
  AOI21X1TF U526 ( .A0(N507), .A1(N331), .B0(N488), .Y(N485) );
  NOR2X1TF U527 ( .A(N314), .B(N480), .Y(N486) );
  INVX2TF U528 ( .A(N501), .Y(N498) );
  AND2X2TF U529 ( .A(\SCPU_CTRL_SPI_FOUT[12] ), .B(N311), .Y(
        \SCPU_CTRL_SPI_IO_DATAINA[12] ) );
  AND2X2TF U530 ( .A(\SCPU_CTRL_SPI_FOUT[11] ), .B(N311), .Y(
        \SCPU_CTRL_SPI_IO_DATAINA[11] ) );
  AOI22X1TF U531 ( .A0(SCPU_CTRL_SPI_D_ADDR[3]), .A1(N404), .B0(N393), .B1(
        N325), .Y(N394) );
  AOI22X1TF U532 ( .A0(Q_FROM_SRAM[2]), .A1(N403), .B0(N402), .B1(
        SCPU_CTRL_SPI_I_ADDR[3]), .Y(N395) );
  AOI22X1TF U533 ( .A0(N401), .A1(\SCPU_CTRL_SPI_IO_DATAINA[2] ), .B0(N400), 
        .B1(\SCPU_CTRL_SPI_POUT[2] ), .Y(N396) );
  AOI22X1TF U534 ( .A0(N399), .A1(I_APP_DONE), .B0(N398), .B1(
        \SCPU_CTRL_SPI_FOUT[2] ), .Y(N397) );
  AOI21X1TF U535 ( .A0(SCPU_CTRL_SPI_D_ADDR[2]), .A1(N404), .B0(N375), .Y(N376) );
  AOI22X1TF U536 ( .A0(N403), .A1(Q_FROM_SRAM[1]), .B0(N402), .B1(
        SCPU_CTRL_SPI_I_ADDR[2]), .Y(N377) );
  AOI22X1TF U537 ( .A0(N401), .A1(\SCPU_CTRL_SPI_IO_DATAINA[1] ), .B0(N400), 
        .B1(\SCPU_CTRL_SPI_POUT[1] ), .Y(N378) );
  AOI22X1TF U538 ( .A0(N399), .A1(N266), .B0(N398), .B1(
        \SCPU_CTRL_SPI_FOUT[1] ), .Y(N379) );
  NOR3X1TF U539 ( .A(N108), .B(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .C(N110), 
        .Y(N266) );
  AOI22X1TF U540 ( .A0(N402), .A1(SCPU_CTRL_SPI_I_ADDR[6]), .B0(N405), .B1(
        SCPU_CTRL_SPI_I_NXT[1]), .Y(N385) );
  AOI22X1TF U541 ( .A0(N400), .A1(\SCPU_CTRL_SPI_POUT[5] ), .B0(N403), .B1(
        Q_FROM_SRAM[5]), .Y(N386) );
  AOI22X1TF U542 ( .A0(N398), .A1(\SCPU_CTRL_SPI_FOUT[5] ), .B0(N401), .B1(
        \SCPU_CTRL_SPI_IO_DATAINA[5] ), .Y(N387) );
  AOI22X1TF U543 ( .A0(N402), .A1(SCPU_CTRL_SPI_I_ADDR[5]), .B0(N405), .B1(
        SCPU_CTRL_SPI_I_NXT[0]), .Y(N381) );
  AOI22X1TF U544 ( .A0(N400), .A1(\SCPU_CTRL_SPI_POUT[4] ), .B0(N403), .B1(
        Q_FROM_SRAM[4]), .Y(N382) );
  AOI22X1TF U545 ( .A0(N398), .A1(\SCPU_CTRL_SPI_FOUT[4] ), .B0(N401), .B1(
        \SCPU_CTRL_SPI_IO_DATAINA[4] ), .Y(N383) );
  AND2X2TF U546 ( .A(\SCPU_CTRL_SPI_FOUT[10] ), .B(N311), .Y(
        \SCPU_CTRL_SPI_IO_DATAINA[10] ) );
  AND3X2TF U547 ( .A(N342), .B(\SCPU_CTRL_SPI_PUT_CNT_STATE[0] ), .C(N405), 
        .Y(N393) );
  AOI22X1TF U548 ( .A0(N403), .A1(Q_FROM_SRAM[3]), .B0(N402), .B1(
        SCPU_CTRL_SPI_I_ADDR[4]), .Y(N390) );
  AOI22X1TF U549 ( .A0(N400), .A1(\SCPU_CTRL_SPI_POUT[3] ), .B0(N404), .B1(
        SCPU_CTRL_SPI_D_ADDR[4]), .Y(N391) );
  AOI22X1TF U550 ( .A0(N398), .A1(\SCPU_CTRL_SPI_FOUT[3] ), .B0(N401), .B1(
        \SCPU_CTRL_SPI_IO_DATAINA[3] ), .Y(N392) );
  AOI22X1TF U551 ( .A0(N405), .A1(SCPU_CTRL_SPI_I_SPI_SO), .B0(N404), .B1(
        SCPU_CTRL_SPI_D_ADDR[1]), .Y(N406) );
  NOR3X2TF U552 ( .A(N374), .B(N373), .C(N372), .Y(N404) );
  INVX2TF U553 ( .A(N388), .Y(N405) );
  AOI22X1TF U554 ( .A0(N403), .A1(Q_FROM_SRAM[0]), .B0(N402), .B1(
        SCPU_CTRL_SPI_I_ADDR[1]), .Y(N407) );
  AOI22X1TF U555 ( .A0(N401), .A1(\SCPU_CTRL_SPI_IO_DATAINA[0] ), .B0(N400), 
        .B1(\SCPU_CTRL_SPI_POUT[0] ), .Y(N408) );
  NOR3X2TF U556 ( .A(I_TEST_MUX[2]), .B(N373), .C(N374), .Y(N400) );
  NOR3X2TF U557 ( .A(I_TEST_MUX[0]), .B(I_TEST_MUX[2]), .C(N374), .Y(N401) );
  AOI22X1TF U558 ( .A0(N399), .A1(\SCPU_CTRL_SPI_IO_STATUS[0] ), .B0(N398), 
        .B1(\SCPU_CTRL_SPI_FOUT[0] ), .Y(N409) );
  NOR3X2TF U559 ( .A(I_TEST_MUX[1]), .B(I_TEST_MUX[2]), .C(N373), .Y(N398) );
  NOR3X1TF U560 ( .A(I_TEST_MUX[1]), .B(I_TEST_MUX[0]), .C(N372), .Y(N399) );
  INVX2TF U561 ( .A(N311), .Y(N474) );
  INVX2TF U562 ( .A(Q_FROM_SRAM[1]), .Y(N466) );
  INVX2TF U563 ( .A(Q_FROM_SRAM[0]), .Y(N465) );
  INVX2TF U564 ( .A(Q_FROM_SRAM[4]), .Y(N469) );
  INVX2TF U565 ( .A(Q_FROM_SRAM[7]), .Y(N473) );
  INVX2TF U566 ( .A(Q_FROM_SRAM[5]), .Y(N470) );
  INVX2TF U567 ( .A(Q_FROM_SRAM[2]), .Y(N467) );
  INVX2TF U568 ( .A(Q_FROM_SRAM[6]), .Y(N471) );
  INVX2TF U569 ( .A(Q_FROM_SRAM[3]), .Y(N468) );
  NAND2X1TF U570 ( .A(N316), .B(N479), .Y(N509) );
  AO21X1TF U571 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ), .A1(N349), .B0(
        N350), .Y(SCPU_CTRL_SPI_CCT_N56) );
  XOR2X1TF U572 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[7] ), .B(N350), .Y(
        SCPU_CTRL_SPI_CCT_N57) );
  AO22X1TF U573 ( .A0(N370), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[1] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[1]), .B1(N439), .Y(D_AFTER_MUX[1]) );
  AO22X1TF U574 ( .A0(N370), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[2] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[2]), .B1(N320), .Y(D_AFTER_MUX[2]) );
  AO22X1TF U575 ( .A0(N370), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[3] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[3]), .B1(N320), .Y(D_AFTER_MUX[3]) );
  AO22X1TF U576 ( .A0(N370), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[4] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[4]), .B1(N320), .Y(D_AFTER_MUX[4]) );
  AO22X1TF U577 ( .A0(N370), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[5] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[5]), .B1(N320), .Y(D_AFTER_MUX[5]) );
  AO22X1TF U578 ( .A0(N370), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[6] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[6]), .B1(N320), .Y(D_AFTER_MUX[6]) );
  AO22X1TF U579 ( .A0(N370), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[7] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[7]), .B1(N320), .Y(D_AFTER_MUX[7]) );
  AO22X1TF U580 ( .A0(N318), .A1(\SCPU_CTRL_SPI_FOUT[1] ), .B0(N474), .B1(
        I_ADC_PI[1]), .Y(\SCPU_CTRL_SPI_IO_DATAINA[1] ) );
  NAND2X1TF U581 ( .A(I_TEST_MUX[0]), .B(I_TEST_MUX[2]), .Y(N371) );
  NAND3X1TF U582 ( .A(N374), .B(N373), .C(N372), .Y(N388) );
  NOR4XLTF U583 ( .A(N110), .B(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .C(N330), 
        .D(N388), .Y(N375) );
  AO22X1TF U584 ( .A0(N311), .A1(\SCPU_CTRL_SPI_FOUT[4] ), .B0(N474), .B1(
        I_ADC_PI[4]), .Y(\SCPU_CTRL_SPI_IO_DATAINA[4] ) );
  NAND2X1TF U585 ( .A(N404), .B(SCPU_CTRL_SPI_D_ADDR[5]), .Y(N380) );
  AO22X1TF U586 ( .A0(N311), .A1(\SCPU_CTRL_SPI_FOUT[5] ), .B0(N474), .B1(
        I_ADC_PI[5]), .Y(\SCPU_CTRL_SPI_IO_DATAINA[5] ) );
  NAND2X1TF U587 ( .A(N404), .B(SCPU_CTRL_SPI_D_ADDR[6]), .Y(N384) );
  AO22X1TF U588 ( .A0(N318), .A1(\SCPU_CTRL_SPI_FOUT[3] ), .B0(N474), .B1(
        I_ADC_PI[3]), .Y(\SCPU_CTRL_SPI_IO_DATAINA[3] ) );
  NAND2X1TF U589 ( .A(\SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .B(N393), .Y(N389) );
  AO22X1TF U590 ( .A0(N311), .A1(\SCPU_CTRL_SPI_FOUT[2] ), .B0(N474), .B1(
        I_ADC_PI[2]), .Y(\SCPU_CTRL_SPI_IO_DATAINA[2] ) );
  AO22X1TF U591 ( .A0(N311), .A1(\SCPU_CTRL_SPI_FOUT[0] ), .B0(N474), .B1(
        I_ADC_PI[0]), .Y(\SCPU_CTRL_SPI_IO_DATAINA[0] ) );
  NAND2BX1TF U592 ( .AN(N264), .B(I_CTRL_MODE[1]), .Y(N263) );
  OAI221XLTF U593 ( .A0(N319), .A1(I_LOAD_N), .B0(N341), .B1(N413), .C0(
        I_CTRL_BGN), .Y(N410) );
  AO22X1TF U594 ( .A0(N319), .A1(N168), .B0(N414), .B1(N410), .Y(N261) );
  NAND2BX1TF U595 ( .AN(I_CTRL_MODE[0]), .B(N416), .Y(N419) );
  NAND2X1TF U596 ( .A(I_CTRL_MODE[0]), .B(N416), .Y(N417) );
  NAND2X1TF U597 ( .A(N108), .B(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .Y(N423) );
  NAND3X1TF U598 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .B(N108), .C(N323), 
        .Y(N442) );
  AOI2BB2X1TF U599 ( .B0(N427), .B1(N323), .A0N(N330), .A1N(
        \SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .Y(N430) );
  NAND2X1TF U600 ( .A(N431), .B(N438), .Y(N433) );
  NAND3X1TF U601 ( .A(N437), .B(N434), .C(N433), .Y(N251) );
  NAND2X1TF U602 ( .A(N438), .B(N334), .Y(N436) );
  OAI2BB2XLTF U603 ( .B0(N473), .B1(N452), .A0N(N450), .A1N(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[7]), .Y(N248) );
  AO22X1TF U604 ( .A0(N311), .A1(\SCPU_CTRL_SPI_FOUT[6] ), .B0(N474), .B1(
        I_ADC_PI[6]), .Y(\SCPU_CTRL_SPI_IO_DATAINA[6] ) );
  AO22X1TF U605 ( .A0(N318), .A1(\SCPU_CTRL_SPI_FOUT[7] ), .B0(N474), .B1(
        I_ADC_PI[7]), .Y(\SCPU_CTRL_SPI_IO_DATAINA[7] ) );
  AO22X1TF U606 ( .A0(N311), .A1(\SCPU_CTRL_SPI_FOUT[8] ), .B0(N474), .B1(
        I_ADC_PI[8]), .Y(\SCPU_CTRL_SPI_IO_DATAINA[8] ) );
  AO22X1TF U607 ( .A0(N318), .A1(\SCPU_CTRL_SPI_FOUT[9] ), .B0(N474), .B1(
        I_ADC_PI[9]), .Y(\SCPU_CTRL_SPI_IO_DATAINA[9] ) );
  AO22X1TF U608 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .A1(
        \SCPU_CTRL_SPI_PUT_CNT_STATE[0] ), .B0(N325), .B1(
        SCPU_CTRL_SPI_PUT_N110), .Y(SCPU_CTRL_SPI_PUT_N111) );
  NAND2X1TF U609 ( .A(N325), .B(N336), .Y(N476) );
  NAND3X1TF U610 ( .A(N328), .B(N324), .C(N515), .Y(N510) );
  NAND3X1TF U611 ( .A(SCPU_CTRL_SPI_A_SPI[2]), .B(SCPU_CTRL_SPI_A_SPI[0]), .C(
        SCPU_CTRL_SPI_A_SPI[1]), .Y(N501) );
  NAND2X1TF U612 ( .A(N498), .B(SCPU_CTRL_SPI_A_SPI[3]), .Y(N497) );
  NOR2BX1TF U613 ( .AN(SCPU_CTRL_SPI_A_SPI[4]), .B(N497), .Y(N491) );
  NAND3X1TF U614 ( .A(N491), .B(SCPU_CTRL_SPI_A_SPI[5]), .C(
        SCPU_CTRL_SPI_A_SPI[6]), .Y(N480) );
  NAND2X1TF U615 ( .A(SCPU_CTRL_SPI_A_SPI[7]), .B(N486), .Y(N483) );
  OAI2BB1X1TF U616 ( .A0N(N480), .A1N(N507), .B0(N509), .Y(N488) );
  AOI2BB2X1TF U617 ( .B0(\SCPU_CTRL_SPI_IO_DATAOUTA[8] ), .B1(N346), .A0N(
        SCPU_CTRL_SPI_A_SPI[8]), .A1N(N483), .Y(N484) );
  OAI2BB1X1TF U618 ( .A0N(SCPU_CTRL_SPI_A_SPI[7]), .A1N(N488), .B0(N487), .Y(
        N94) );
  NAND2X1TF U619 ( .A(N507), .B(N491), .Y(N494) );
  XNOR2X1TF U621 ( .A(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .B(N512), .Y(N36)
         );
endmodule

