
module SHARE_SUPERALU_VG ( CLK, RST_N, X_IN, Y_IN, ALU_START, ALU_TYPE, MODE_TYPE, 
        OFFSET, FOUT, POUT, ALU_IS_DONE );
  input [12:0] X_IN;
  input [12:0] Y_IN;
  input [2:0] ALU_TYPE;
  input [1:0] MODE_TYPE;
  input [9:0] OFFSET;
  output [12:0] FOUT;
  output [12:0] POUT;
  input CLK, RST_N, ALU_START;
  output ALU_IS_DONE;
  wire   POST_WORK, PRE_WORK, \INDEX[2] , \RSHT_BITS[3] , SIGN_Y, C152_DATA4_0,
         C152_DATA4_1, C152_DATA4_2, C152_DATA4_3, C152_DATA4_4, C152_DATA4_5,
         C152_DATA4_6, C152_DATA4_7, C152_DATA4_8, C152_DATA4_9, C152_DATA4_10,
         C152_DATA4_11, C152_DATA4_12, N74, N90, N91, N92, N121, N122, N123,
         N124, N128, N129, N657, N658, N659, N660, N661, N662, N663, N664,
         N665, N666, N667, N668, N669, N670, N671, N672, N673, N674, N675,
         N676, N677, N678, N679, N680, N681, N682, N683, N684, N685, N686,
         N687, N688, N689, N690, N691, N692, N693, N694, N695, N696, N697,
         N698, N699, N700, N701, N702, N703, N704, N705, N706, N707, N708,
         N709, N710, N711, N712, N713, N714, N715, N716, N717, N718, N719,
         N720, N721, N722, N723, N724, N725, N726, C2_Z_12, C2_Z_11, C2_Z_10,
         C2_Z_9, C2_Z_8, C2_Z_7, C2_Z_5, C2_Z_4, C2_Z_3, C2_Z_2, C2_Z_1,
         INTADD_0_CI, \INTADD_0_SUM[6] , \INTADD_0_SUM[5] , \INTADD_0_SUM[4] ,
         \INTADD_0_SUM[3] , \INTADD_0_SUM[2] , \INTADD_0_SUM[1] ,
         \INTADD_0_SUM[0] , INTADD_0_N7, INTADD_0_N6, INTADD_0_N5, INTADD_0_N4,
         INTADD_0_N3, INTADD_0_N2, INTADD_0_N1, ADD_X_132_1_N13,
         ADD_X_132_1_N12, ADD_X_132_1_N11, ADD_X_132_1_N10, ADD_X_132_1_N9,
         ADD_X_132_1_N8, ADD_X_132_1_N7, ADD_X_132_1_N6, ADD_X_132_1_N5,
         ADD_X_132_1_N4, ADD_X_132_1_N3, ADD_X_132_1_N2,
         DP_OP_333_124_4748_N57, DP_OP_333_124_4748_N43,
         DP_OP_333_124_4748_N28, DP_OP_333_124_4748_N27,
         DP_OP_333_124_4748_N26, DP_OP_333_124_4748_N25,
         DP_OP_333_124_4748_N24, DP_OP_333_124_4748_N22,
         DP_OP_333_124_4748_N21, DP_OP_333_124_4748_N20,
         DP_OP_333_124_4748_N19, DP_OP_333_124_4748_N18,
         DP_OP_333_124_4748_N17, DP_OP_333_124_4748_N12,
         DP_OP_333_124_4748_N11, DP_OP_333_124_4748_N10, DP_OP_333_124_4748_N9,
         DP_OP_333_124_4748_N8, DP_OP_333_124_4748_N7, DP_OP_333_124_4748_N6,
         DP_OP_333_124_4748_N5, DP_OP_333_124_4748_N4, DP_OP_333_124_4748_N3,
         DP_OP_333_124_4748_N2, DP_OP_333_124_4748_N1, N1, N2, N3, N4, N5, N6,
         N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62,
         N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N75, N76, N77,
         N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N93, N94,
         N95, N96, N97, N98, N99, N100, N119, N120, N125, N126, N127, N130,
         N131, N132, N133, N134, N135, N136, N137, N138, N139, N140, N141,
         N142, N143, N144, N145, N146, N147, N148, N149, N150, N151, N152,
         N153, N154, N155, N156, N157, N158, N159, N160, N161, N162, N163,
         N164, N165, N166, N167, N168, N169, N170, N171, N172, N173, N174,
         N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N185,
         N186, N187, N188, N189, N190, N191, N192, N193, N194, N195, N196,
         N197, N198, N199, N200, N201, N202, N203, N204, N205, N206, N207,
         N208, N209, N210, N211, N212, N213, N214, N215, N216, N217, N218,
         N219, N220, N221, N222, N223, N224, N225, N226, N227, N228, N229,
         N230, N231, N232, N233, N234, N235, N236, N237, N238, N239, N240,
         N241, N242, N243, N244, N245, N246, N247, N248, N249, N250, N251,
         N252, N253, N254, N255, N256, N257, N258, N259, N260, N261, N262,
         N263, N264, N265, N266, N267, N268, N269, N270, N271, N272, N273,
         N274, N275, N276, N277, N278, N279, N280, N281, N282, N283, N284,
         N285, N286, N287, N288, N289, N290, N291, N292, N293, N294, N295,
         N296, N297, N298, N299, N300, N301, N302, N303, N304, N305, N306,
         N307, N308, N309, N310, N311, N312, N313, N314, N315, N316, N317,
         N318, N319, N320, N321, N322, N323, N324, N325, N326, N327, N328,
         N329, N330, N331, N332, N333, N334, N335, N336, N337, N338, N339,
         N340, N341, N342, N343, N344, N345, N346, N347, N348, N349, N350,
         N351, N352, N353, N354, N355, N356, N357, N358, N359, N360, N361,
         N362, N363, N364, N365, N366, N367, N368, N369, N370, N371, N372,
         N373, N374, N375, N376, N377, N378, N379, N380, N381, N382, N383,
         N384, N385, N386, N387, N388, N389, N390, N391, N392, N393, N394,
         N395, N396, N397, N398, N399, N400, N401, N402, N403, N404, N405,
         N406, N407, N408, N409, N410, N411, N412, N413, N414, N415, N416,
         N417, N418, N419, N420, N421, N422, N423, N424, N425, N426, N427,
         N428, N429, N430, N431, N432, N433, N434, N435, N436, N437, N438,
         N439, N440, N441, N442, N443, N444, N445, N446, N447, N448, N449,
         N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460,
         N461, N462, N463, N464, N465, N466, N467, N468, N469, N470, N471,
         N472, N473, N474, N475, N476, N477, N478, N479, N480, N481, N482,
         N483, N484, N485, N486, N487, N488, N489, N490, N491, N492, N493,
         N494, N495, N496, N497, N498, N499, N500, N501, N502, N503, N504,
         N505, N506, N507, N508, N509, N510, N511, N512, N513, N514, N515,
         N516, N517, N518, N519, N520, N521, N522, N523, N524, N525, N526,
         N527, N528, N529, N530, N531, N532, N533, N534, N535, N536, N537,
         N538, N539, N540, N541, N542, N543, N544, N545, N546, N547, N548,
         N549, N550, N551, N552, N553, N554, N555, N556, N557, N558, N559,
         N560, N561, N562, N563, N564, N565, N566, N567, N568, N569, N570,
         N571, N572, N573, N574, N575, N576, N577, N578, N579, N580, N581,
         N582, N583, N584, N585, N586, N587, N588, N589, N590, N591, N592,
         N593, N594, N595, N596, N597, N598, N599, N600, N601, N602, N603,
         N604, N605, N606, N607, N608, N609, N610, N611, N612, N613, N614,
         N615, N616, N617, N618, N619, N620, N621, N622, N623, N624, N625,
         N626, N627, N628, N629, N630, N631, N632, N633, N634, N635, N636,
         N637, N638, N639, N640, N641, N642, N643, N644, N645, N646, N647,
         N648, N649, N650, N651, N652, N653, N654, N655, N656, N727, N728,
         N729, N730, N731, N732, N733, N734, N735, N736, N737, N738, N739,
         N740, N741, N742, N743, N744, N745, N746, N747, N748, N749, N750,
         N751, N752, N753, N754, N755, N756, N757, N758, N759, N760, N761,
         N762, N763, N764, N765, N766, N767, N768, N769, N770, N771, N772,
         N773, N774, N775, N776, N777, N778, N779, N780, N781, N782, N783,
         N784, N785, N786, N787, N788, N789, N790, N791, N792, N793, N794,
         N795, N796, N797, N798, N799, N800, N801, N802, N803, N804, N805,
         N806, N807, N808, N809, N810, N811, N812, N813, N814, N815, N816,
         N817, N818, N819, N820, N821, N822, N823, N824, N825, N826, N827,
         N828, N829, N830, N831, N832, N833, N834, N835, N836, N837, N838,
         N839, N840, N841, N842, N843, N844, N845, N846, N847, N848, N849,
         N850, N851, N852, N853, N854, N855, N856, N857, N858, N859, N860,
         N861, N862, N863, N864, N865, N866, N867, N868, N869, N870, N871,
         N872, N873, N874, N875, N876, N877, N878, N879, N880, N881, N882,
         N883, N884, N885, N886, N887, N888, N889, N890, N891, N892, N893,
         N894, N895, N896, N897, N898, N899, N900, N901, N902, N903, N904,
         N905, N906, N907, N908, N909, N910, N911, N912, N913, N914, N915,
         N916, N917, N918, N919, N920, N921, N922, N923, N924, N925, N926,
         N927, N928, N929, N930, N931, N932, N933, N934, N935, N936, N937,
         N938, N939, N940, N941, N942, N943, N944, N945, N946, N947, N948,
         N949, N950, N951, N952, N953, N954, N955, N956, N957, N958, N959,
         N960, N961, N962, N963, N964, N965, N966, N967, N968, N969, N970,
         N971, N972, N973, N974, N975, N976, N977, N978, N979, N980, N981,
         N982, N983, N984, N985, N986, N987, N988, N989, N990, N991, N992,
         N993, N994, N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003,
         N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013,
         N1014, N1015, N1016, N1017, N1018;
  wire   [12:9] XTEMP;
  wire   [12:0] DIVISION_HEAD;
  wire   [8:0] DIVISION_REMA;
  wire   [12:0] OPER_A;
  wire   [12:0] OPER_B;
  wire   [12:0] SUM_AB;
  wire   [12:0] ZTEMP;
  wire   [3:2] STEP;

  CMPR32X2TF \intadd_0/U7  ( .A(N174), .B(DIVISION_HEAD[6]), .C(INTADD_0_N7), 
        .CO(INTADD_0_N6), .S(\INTADD_0_SUM[1] ) );
  CMPR32X2TF \intadd_0/U6  ( .A(N56), .B(DIVISION_HEAD[7]), .C(INTADD_0_N6), 
        .CO(INTADD_0_N5), .S(\INTADD_0_SUM[2] ) );
  CMPR32X2TF \intadd_0/U5  ( .A(N175), .B(DIVISION_HEAD[8]), .C(INTADD_0_N5), 
        .CO(INTADD_0_N4), .S(\INTADD_0_SUM[3] ) );
  CMPR32X2TF \intadd_0/U4  ( .A(N61), .B(DIVISION_HEAD[9]), .C(INTADD_0_N4), 
        .CO(INTADD_0_N3), .S(\INTADD_0_SUM[4] ) );
  CMPR32X2TF \intadd_0/U3  ( .A(X_IN[6]), .B(DIVISION_HEAD[10]), .C(
        INTADD_0_N3), .CO(INTADD_0_N2), .S(\INTADD_0_SUM[5] ) );
  CMPR32X2TF \intadd_0/U2  ( .A(N176), .B(DIVISION_HEAD[11]), .C(INTADD_0_N2), 
        .CO(INTADD_0_N1), .S(\INTADD_0_SUM[6] ) );
  DFFRX2TF \wtemp_reg[9]  ( .D(N673), .CK(CLK), .RN(RST_N), .Q(OPER_B[9]), 
        .QN(N168) );
  DFFRX2TF \wtemp_reg[12]  ( .D(N724), .CK(CLK), .RN(RST_N), .Q(OPER_B[12]), 
        .QN(N167) );
  DFFRX2TF \index_reg[3]  ( .D(N725), .CK(CLK), .RN(RST_N), .Q(N166), .QN(N124) );
  DFFRX2TF \wtemp_reg[11]  ( .D(N671), .CK(CLK), .RN(RST_N), .Q(OPER_B[11]), 
        .QN(N165) );
  DFFRX2TF \wtemp_reg[0]  ( .D(N682), .CK(CLK), .RN(RST_N), .Q(OPER_B[0]), 
        .QN(N164) );
  DFFSX2TF pre_work_reg ( .D(N695), .CK(CLK), .SN(RST_N), .Q(PRE_WORK), .QN(
        N156) );
  DFFRX2TF \wtemp_reg[4]  ( .D(N678), .CK(CLK), .RN(RST_N), .Q(OPER_B[4]), 
        .QN(N155) );
  DFFRX2TF \ytemp_reg[10]  ( .D(N684), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[1]), .QN(N150) );
  DFFRX2TF \ytemp_reg[9]  ( .D(N685), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[0]), .QN(N148) );
  DFFRX2TF \ytemp_reg[8]  ( .D(N686), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[8]), .QN(N144) );
  DFFRX2TF \xtemp_reg[10]  ( .D(N709), .CK(CLK), .RN(RST_N), .Q(XTEMP[10]), 
        .QN(N136) );
  DFFRX2TF \xtemp_reg[11]  ( .D(N708), .CK(CLK), .RN(RST_N), .Q(XTEMP[11]), 
        .QN(N133) );
  DFFRX2TF \xtemp_reg[0]  ( .D(N719), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[4]), .QN(N125) );
  DFFRX2TF \rsht_bits_reg[2]  ( .D(N701), .CK(CLK), .RN(RST_N), .QN(N90) );
  DFFRX2TF \index_reg[2]  ( .D(N698), .CK(CLK), .RN(RST_N), .Q(\INDEX[2] ) );
  DFFRX2TF \ztemp_reg[12]  ( .D(N657), .CK(CLK), .RN(RST_N), .Q(ZTEMP[12]) );
  DFFRX2TF \ztemp_reg[11]  ( .D(N658), .CK(CLK), .RN(RST_N), .Q(ZTEMP[11]) );
  DFFRX2TF \ztemp_reg[10]  ( .D(N659), .CK(CLK), .RN(RST_N), .Q(ZTEMP[10]) );
  DFFRX2TF \ztemp_reg[9]  ( .D(N660), .CK(CLK), .RN(RST_N), .Q(ZTEMP[9]) );
  DFFRX2TF \wtemp_reg[6]  ( .D(N676), .CK(CLK), .RN(RST_N), .Q(OPER_B[6]) );
  DFFRX2TF \wtemp_reg[7]  ( .D(N675), .CK(CLK), .RN(RST_N), .Q(OPER_B[7]) );
  DFFRX2TF \ztemp_reg[8]  ( .D(N661), .CK(CLK), .RN(RST_N), .Q(ZTEMP[8]) );
  DFFRX2TF \ztemp_reg[7]  ( .D(N662), .CK(CLK), .RN(RST_N), .Q(ZTEMP[7]) );
  DFFRX2TF \ztemp_reg[6]  ( .D(N663), .CK(CLK), .RN(RST_N), .Q(ZTEMP[6]) );
  DFFRX2TF \ztemp_reg[5]  ( .D(N664), .CK(CLK), .RN(RST_N), .Q(ZTEMP[5]) );
  DFFRX2TF \ztemp_reg[4]  ( .D(N665), .CK(CLK), .RN(RST_N), .Q(ZTEMP[4]) );
  DFFRX2TF \xtemp_reg[9]  ( .D(N710), .CK(CLK), .RN(RST_N), .Q(XTEMP[9]), .QN(
        N39) );
  DFFRX2TF \wtemp_reg[5]  ( .D(N677), .CK(CLK), .RN(RST_N), .Q(OPER_B[5]) );
  DFFRX2TF \ytemp_reg[12]  ( .D(N706), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[3]), .QN(N40) );
  DFFRX2TF \ytemp_reg[11]  ( .D(N683), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[2]), .QN(N43) );
  DFFRX2TF \xtemp_reg[12]  ( .D(N723), .CK(CLK), .RN(RST_N), .Q(XTEMP[12]), 
        .QN(N44) );
  DFFRX2TF \ztemp_reg[3]  ( .D(N666), .CK(CLK), .RN(RST_N), .Q(ZTEMP[3]) );
  DFFRX2TF \ztemp_reg[2]  ( .D(N667), .CK(CLK), .RN(RST_N), .Q(ZTEMP[2]) );
  DFFRX2TF \ztemp_reg[1]  ( .D(N668), .CK(CLK), .RN(RST_N), .Q(ZTEMP[1]) );
  DFFRX2TF \ztemp_reg[0]  ( .D(N669), .CK(CLK), .RN(RST_N), .Q(ZTEMP[0]) );
  DFFRX2TF \xtemp_reg[3]  ( .D(N716), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[7]), .QN(N42) );
  CMPR32X2TF \add_x_132_1/U4  ( .A(OPER_A[10]), .B(OPER_B[10]), .C(
        ADD_X_132_1_N4), .CO(ADD_X_132_1_N3), .S(SUM_AB[10]) );
  CMPR32X2TF \add_x_132_1/U8  ( .A(OPER_A[6]), .B(OPER_B[6]), .C(
        ADD_X_132_1_N8), .CO(ADD_X_132_1_N7), .S(SUM_AB[6]) );
  CMPR32X2TF \add_x_132_1/U10  ( .A(OPER_A[4]), .B(OPER_B[4]), .C(
        ADD_X_132_1_N10), .CO(ADD_X_132_1_N9), .S(SUM_AB[4]) );
  CMPR32X2TF \add_x_132_1/U13  ( .A(OPER_A[1]), .B(OPER_B[1]), .C(
        ADD_X_132_1_N13), .CO(ADD_X_132_1_N12), .S(SUM_AB[1]) );
  CMPR32X2TF \add_x_132_1/U5  ( .A(OPER_A[9]), .B(OPER_B[9]), .C(
        ADD_X_132_1_N5), .CO(ADD_X_132_1_N4), .S(SUM_AB[9]) );
  CMPR32X2TF \add_x_132_1/U12  ( .A(OPER_A[2]), .B(OPER_B[2]), .C(
        ADD_X_132_1_N12), .CO(ADD_X_132_1_N11), .S(SUM_AB[2]) );
  CMPR32X2TF \add_x_132_1/U11  ( .A(OPER_A[3]), .B(OPER_B[3]), .C(
        ADD_X_132_1_N11), .CO(ADD_X_132_1_N10), .S(SUM_AB[3]) );
  CMPR32X2TF \add_x_132_1/U9  ( .A(OPER_A[5]), .B(OPER_B[5]), .C(
        ADD_X_132_1_N9), .CO(ADD_X_132_1_N8), .S(SUM_AB[5]) );
  CMPR32X2TF \add_x_132_1/U7  ( .A(OPER_A[7]), .B(OPER_B[7]), .C(
        ADD_X_132_1_N7), .CO(ADD_X_132_1_N6), .S(SUM_AB[7]) );
  CMPR32X2TF \add_x_132_1/U3  ( .A(OPER_A[11]), .B(OPER_B[11]), .C(
        ADD_X_132_1_N3), .CO(ADD_X_132_1_N2), .S(SUM_AB[11]) );
  ADDHX1TF \DP_OP_333_124_4748/U5  ( .A(DP_OP_333_124_4748_N21), .B(
        DP_OP_333_124_4748_N5), .CO(DP_OP_333_124_4748_N4), .S(C152_DATA4_8)
         );
  ADDHXLTF \DP_OP_333_124_4748/U11  ( .A(DP_OP_333_124_4748_N27), .B(
        DP_OP_333_124_4748_N11), .CO(DP_OP_333_124_4748_N10), .S(C152_DATA4_2)
         );
  ADDHXLTF \DP_OP_333_124_4748/U10  ( .A(DP_OP_333_124_4748_N26), .B(
        DP_OP_333_124_4748_N10), .CO(DP_OP_333_124_4748_N9), .S(C152_DATA4_3)
         );
  ADDHX1TF \DP_OP_333_124_4748/U6  ( .A(DP_OP_333_124_4748_N22), .B(
        DP_OP_333_124_4748_N6), .CO(DP_OP_333_124_4748_N5), .S(C152_DATA4_7)
         );
  ADDHXLTF \DP_OP_333_124_4748/U12  ( .A(DP_OP_333_124_4748_N28), .B(
        DP_OP_333_124_4748_N12), .CO(DP_OP_333_124_4748_N11), .S(C152_DATA4_1)
         );
  ADDHX1TF \DP_OP_333_124_4748/U2  ( .A(DP_OP_333_124_4748_N18), .B(
        DP_OP_333_124_4748_N2), .CO(DP_OP_333_124_4748_N1), .S(C152_DATA4_11)
         );
  ADDHX1TF \DP_OP_333_124_4748/U4  ( .A(DP_OP_333_124_4748_N20), .B(
        DP_OP_333_124_4748_N4), .CO(DP_OP_333_124_4748_N3), .S(C152_DATA4_9)
         );
  ADDHX1TF \DP_OP_333_124_4748/U3  ( .A(DP_OP_333_124_4748_N19), .B(
        DP_OP_333_124_4748_N3), .CO(DP_OP_333_124_4748_N2), .S(C152_DATA4_10)
         );
  XOR2X1TF \DP_OP_333_124_4748/U27  ( .A(DP_OP_333_124_4748_N43), .B(C2_Z_1), 
        .Y(DP_OP_333_124_4748_N28) );
  XOR2X1TF \DP_OP_333_124_4748/U26  ( .A(DP_OP_333_124_4748_N43), .B(C2_Z_2), 
        .Y(DP_OP_333_124_4748_N27) );
  XOR2X1TF \DP_OP_333_124_4748/U25  ( .A(N93), .B(C2_Z_3), .Y(
        DP_OP_333_124_4748_N26) );
  XOR2X1TF \DP_OP_333_124_4748/U24  ( .A(N93), .B(C2_Z_4), .Y(
        DP_OP_333_124_4748_N25) );
  XOR2X1TF \DP_OP_333_124_4748/U23  ( .A(N93), .B(C2_Z_5), .Y(
        DP_OP_333_124_4748_N24) );
  XOR2X1TF \DP_OP_333_124_4748/U21  ( .A(N93), .B(C2_Z_7), .Y(
        DP_OP_333_124_4748_N22) );
  XOR2X1TF \DP_OP_333_124_4748/U20  ( .A(N93), .B(C2_Z_8), .Y(
        DP_OP_333_124_4748_N21) );
  XOR2X1TF \DP_OP_333_124_4748/U19  ( .A(N93), .B(C2_Z_9), .Y(
        DP_OP_333_124_4748_N20) );
  XOR2X1TF \DP_OP_333_124_4748/U18  ( .A(N93), .B(C2_Z_10), .Y(
        DP_OP_333_124_4748_N19) );
  XOR2X1TF \DP_OP_333_124_4748/U17  ( .A(N93), .B(C2_Z_11), .Y(
        DP_OP_333_124_4748_N18) );
  XOR2X1TF \DP_OP_333_124_4748/U16  ( .A(N93), .B(C2_Z_12), .Y(
        DP_OP_333_124_4748_N17) );
  XOR2X1TF \DP_OP_333_124_4748/U1  ( .A(DP_OP_333_124_4748_N1), .B(
        DP_OP_333_124_4748_N17), .Y(C152_DATA4_12) );
  DFFRX2TF sign_x_reg ( .D(N722), .CK(CLK), .RN(RST_N), .Q(N963), .QN(N74) );
  DFFRX2TF sign_y_reg ( .D(N694), .CK(CLK), .RN(RST_N), .Q(SIGN_Y), .QN(N157)
         );
  DFFRX2TF XOR_SRC_reg ( .D(N707), .CK(CLK), .RN(RST_N), .Q(N45), .QN(N64) );
  DFFRX2TF SEL_Z_reg ( .D(N670), .CK(CLK), .RN(RST_N), .Q(N142), .QN(N123) );
  DFFRX2TF \step_reg[1]  ( .D(N700), .CK(CLK), .RN(RST_N), .Q(N147), .QN(N121)
         );
  DFFRX2TF \step_reg[2]  ( .D(N696), .CK(CLK), .RN(RST_N), .Q(STEP[2]), .QN(
        N134) );
  DFFRX2TF \step_reg[3]  ( .D(N721), .CK(CLK), .RN(RST_N), .Q(STEP[3]), .QN(
        N149) );
  DFFRX2TF \step_reg[0]  ( .D(N697), .CK(CLK), .RN(RST_N), .Q(N120), .QN(N122)
         );
  DFFRX2TF SEL_SRC_reg ( .D(N720), .CK(CLK), .RN(RST_N), .Q(POST_WORK), .QN(
        N141) );
  DFFRX2TF \rsht_bits_reg[1]  ( .D(N702), .CK(CLK), .RN(RST_N), .Q(N138), .QN(
        N91) );
  DFFRX2TF \rsht_bits_reg[0]  ( .D(N703), .CK(CLK), .RN(RST_N), .Q(N159), .QN(
        N92) );
  DFFRX2TF \index_reg[0]  ( .D(N726), .CK(CLK), .RN(RST_N), .Q(N137), .QN(N129) );
  DFFRX2TF \wtemp_reg[10]  ( .D(N672), .CK(CLK), .RN(RST_N), .Q(OPER_B[10]), 
        .QN(N140) );
  DFFRX2TF \ytemp_reg[1]  ( .D(N693), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[1]), .QN(N158) );
  DFFRX2TF \ytemp_reg[0]  ( .D(N705), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[0]), .QN(N161) );
  DFFRX2TF \rsht_bits_reg[3]  ( .D(N704), .CK(CLK), .RN(RST_N), .Q(
        \RSHT_BITS[3] ), .QN(N169) );
  DFFRX2TF \ytemp_reg[7]  ( .D(N687), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[7]), .QN(N146) );
  DFFRX2TF \wtemp_reg[8]  ( .D(N674), .CK(CLK), .RN(RST_N), .Q(OPER_B[8]), 
        .QN(N139) );
  DFFRX2TF \index_reg[1]  ( .D(N699), .CK(CLK), .RN(RST_N), .Q(N160), .QN(N128) );
  DFFRX2TF \ytemp_reg[6]  ( .D(N688), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[6]), .QN(N152) );
  DFFRX2TF \ytemp_reg[4]  ( .D(N690), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[4]), .QN(N151) );
  DFFRX2TF \ytemp_reg[2]  ( .D(N692), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[2]), .QN(N153) );
  DFFRX2TF \ytemp_reg[5]  ( .D(N689), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[5]), .QN(N145) );
  DFFRX2TF \ytemp_reg[3]  ( .D(N691), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[3]), .QN(N143) );
  DFFRX2TF \xtemp_reg[6]  ( .D(N713), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[10]), .QN(N132) );
  DFFRX2TF \wtemp_reg[2]  ( .D(N680), .CK(CLK), .RN(RST_N), .Q(OPER_B[2]), 
        .QN(N154) );
  DFFRX2TF \xtemp_reg[5]  ( .D(N714), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[9]), .QN(N131) );
  DFFRX2TF \xtemp_reg[2]  ( .D(N717), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[6]), .QN(N126) );
  DFFRX2TF \xtemp_reg[4]  ( .D(N715), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[8]), .QN(N130) );
  DFFRX2TF \wtemp_reg[1]  ( .D(N681), .CK(CLK), .RN(RST_N), .Q(OPER_B[1]), 
        .QN(N162) );
  DFFRX2TF \xtemp_reg[7]  ( .D(N712), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[11]), .QN(N127) );
  DFFRX2TF \xtemp_reg[1]  ( .D(N718), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[5]), .QN(N119) );
  DFFRX2TF \xtemp_reg[8]  ( .D(N711), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[12]), .QN(N135) );
  DFFRX2TF \wtemp_reg[3]  ( .D(N679), .CK(CLK), .RN(RST_N), .Q(OPER_B[3]), 
        .QN(N163) );
  NAND2X2TF U3 ( .A(N307), .B(N655), .Y(N309) );
  INVX2TF U4 ( .A(N243), .Y(N48) );
  NOR2X1TF U5 ( .A(N45), .B(N906), .Y(N895) );
  NAND2X1TF U6 ( .A(X_IN[6]), .B(N729), .Y(N272) );
  NOR2X1TF U7 ( .A(PRE_WORK), .B(N333), .Y(N335) );
  OAI21X2TF U8 ( .A0(X_IN[12]), .A1(N781), .B0(N283), .Y(N767) );
  NAND2X1TF U9 ( .A(N919), .B(N140), .Y(N933) );
  INVX2TF U10 ( .A(N81), .Y(DP_OP_333_124_4748_N43) );
  CLKBUFX2TF U11 ( .A(N244), .Y(N97) );
  NAND2X1TF U12 ( .A(N771), .B(N763), .Y(N396) );
  NOR2X1TF U13 ( .A(OPER_B[1]), .B(OPER_B[0]), .Y(N834) );
  INVX2TF U14 ( .A(N906), .Y(N206) );
  INVX2TF U15 ( .A(N175), .Y(N443) );
  INVX2TF U16 ( .A(Y_IN[0]), .Y(N655) );
  NOR2X1TF U17 ( .A(OPER_A[7]), .B(N879), .Y(N886) );
  NAND2X1TF U18 ( .A(N646), .B(N58), .Y(N946) );
  INVX2TF U19 ( .A(N928), .Y(N931) );
  CLKBUFX2TF U20 ( .A(N734), .Y(N47) );
  NOR2X1TF U21 ( .A(OPER_A[5]), .B(N855), .Y(N865) );
  BUFX3TF U22 ( .A(N49), .Y(N171) );
  NOR2X1TF U23 ( .A(N1017), .B(N1013), .Y(N1012) );
  NAND2X1TF U24 ( .A(N129), .B(N128), .Y(N620) );
  INVX2TF U25 ( .A(N461), .Y(N476) );
  CLKBUFX2TF U26 ( .A(N779), .Y(N170) );
  CLKBUFX6TF U27 ( .A(X_IN[4]), .Y(N175) );
  NOR2X1TF U28 ( .A(OPER_A[3]), .B(N836), .Y(N845) );
  OAI21X2TF U29 ( .A0(N125), .A1(N48), .B0(N229), .Y(OPER_A[0]) );
  NAND2X1TF U30 ( .A(N892), .B(N860), .Y(N882) );
  NOR2X1TF U31 ( .A(\INDEX[2] ), .B(N620), .Y(N305) );
  OR3X1TF U32 ( .A(N871), .B(N870), .C(N196), .Y(N676) );
  OAI22X1TF U33 ( .A0(N185), .A1(OFFSET[4]), .B0(N81), .B1(N180), .Y(N1) );
  XOR2X1TF U34 ( .A(N93), .B(N1), .Y(N2) );
  AND2X2TF U35 ( .A(DP_OP_333_124_4748_N7), .B(N2), .Y(DP_OP_333_124_4748_N6)
         );
  XOR2X1TF U36 ( .A(DP_OP_333_124_4748_N7), .B(N2), .Y(C152_DATA4_6) );
  CLKINVX1TF U37 ( .A(N834), .Y(N3) );
  AOI211X1TF U38 ( .A0(N829), .A1(N830), .B0(N912), .C0(OPER_A[2]), .Y(N4) );
  AOI31X1TF U39 ( .A0(N918), .A1(N154), .A2(N3), .B0(N4), .Y(N5) );
  OAI31X1TF U40 ( .A0(OPER_A[0]), .A1(OPER_A[1]), .A2(N912), .B0(N833), .Y(N6)
         );
  AOI22X1TF U41 ( .A0(OPER_B[3]), .A1(N916), .B0(OPER_A[2]), .B1(N6), .Y(N7)
         );
  AOI32X1TF U42 ( .A0(N918), .A1(OPER_B[2]), .A2(N834), .B0(N917), .B1(
        OPER_B[2]), .Y(N8) );
  AOI31X1TF U43 ( .A0(N5), .A1(N7), .A2(N8), .B0(N920), .Y(N9) );
  AND4X1TF U44 ( .A(N963), .B(N45), .C(N157), .D(N206), .Y(N10) );
  OAI2BB2XLTF U45 ( .B0(N154), .B1(N925), .A0N(N88), .A1N(C152_DATA4_2), .Y(
        N11) );
  OR4X1TF U46 ( .A(N871), .B(N9), .C(N10), .D(N11), .Y(N680) );
  CLKINVX1TF U47 ( .A(N854), .Y(N12) );
  OAI31X1TF U48 ( .A0(OPER_B[5]), .A1(N934), .A2(N12), .B0(N893), .Y(N13) );
  AOI21X1TF U49 ( .A0(C152_DATA4_5), .A1(N88), .B0(N13), .Y(N14) );
  NOR2X1TF U50 ( .A(N931), .B(OPER_A[5]), .Y(N15) );
  AOI22X1TF U51 ( .A0(N855), .A1(N15), .B0(OPER_B[6]), .B1(N853), .Y(N16) );
  OAI21X1TF U52 ( .A0(N854), .A1(N934), .B0(N932), .Y(N17) );
  OAI21X1TF U53 ( .A0(N855), .A1(N931), .B0(N929), .Y(N18) );
  AOI22X1TF U54 ( .A0(OPER_B[5]), .A1(N17), .B0(OPER_A[5]), .B1(N18), .Y(N19)
         );
  NAND4X1TF U55 ( .A(N856), .B(N14), .C(N16), .D(N19), .Y(N677) );
  AOI32X1TF U56 ( .A0(N89), .A1(N835), .A2(N932), .B0(N164), .B1(N835), .Y(N20) );
  AOI211X1TF U57 ( .A0(C152_DATA4_0), .A1(N88), .B0(N874), .C0(N20), .Y(N21)
         );
  OAI21X1TF U58 ( .A0(N844), .A1(N928), .B0(OPER_A[0]), .Y(N22) );
  OAI211X1TF U59 ( .A0(N162), .A1(N882), .B0(N21), .C0(N22), .Y(N682) );
  AOI2BB2X1TF U60 ( .B0(N176), .B1(N274), .A0N(N489), .A1N(N172), .Y(N23) );
  CLKINVX1TF U61 ( .A(Y_IN[4]), .Y(N24) );
  OAI21X1TF U62 ( .A0(N274), .A1(N176), .B0(N24), .Y(N25) );
  AOI22X1TF U63 ( .A0(N489), .A1(N172), .B0(N23), .B1(N25), .Y(N277) );
  AOI21X1TF U64 ( .A0(N200), .A1(C152_DATA4_7), .B0(N189), .Y(N26) );
  OAI31X1TF U65 ( .A0(N875), .A1(N934), .A2(OPER_B[7]), .B0(N26), .Y(N876) );
  OAI21X1TF U66 ( .A0(N82), .A1(N655), .B0(N185), .Y(N27) );
  CLKMX2X2TF U67 ( .A(DP_OP_333_124_4748_N43), .B(DP_OP_333_124_4748_N57), 
        .S0(N27), .Y(DP_OP_333_124_4748_N12) );
  XOR2X1TF U68 ( .A(DP_OP_333_124_4748_N57), .B(N27), .Y(C152_DATA4_0) );
  OAI21X1TF U69 ( .A0(N305), .A1(N628), .B0(N621), .Y(N28) );
  AOI21X1TF U70 ( .A0(N166), .A1(N28), .B0(N383), .Y(N29) );
  NAND4X1TF U71 ( .A(N124), .B(N617), .C(N624), .D(\INDEX[2] ), .Y(N30) );
  NAND4X1TF U72 ( .A(N361), .B(N29), .C(N802), .D(N30), .Y(N725) );
  AOI2BB2X1TF U73 ( .B0(X_IN[6]), .B1(N288), .A0N(Y_IN[5]), .A1N(N469), .Y(N31) );
  CLKINVX1TF U74 ( .A(Y_IN[4]), .Y(N32) );
  OAI21X1TF U75 ( .A0(N288), .A1(X_IN[6]), .B0(N32), .Y(N33) );
  AOI22X1TF U76 ( .A0(N172), .A1(N469), .B0(N31), .B1(N33), .Y(N291) );
  AOI21X1TF U77 ( .A0(N875), .A1(N898), .B0(N873), .Y(N34) );
  NOR2BX1TF U78 ( .AN(OPER_B[7]), .B(N34), .Y(N877) );
  NOR3X1TF U79 ( .A(N950), .B(N949), .C(N81), .Y(N35) );
  AOI211X1TF U80 ( .A0(N944), .A1(N948), .B0(N968), .C0(N35), .Y(N36) );
  OAI22X1TF U81 ( .A0(N943), .A1(N75), .B0(N942), .B1(N971), .Y(N37) );
  NOR4XLTF U82 ( .A(N947), .B(N945), .C(N946), .D(N37), .Y(N38) );
  MXI2X1TF U83 ( .A(N36), .B(N123), .S0(N38), .Y(N670) );
  OAI32X4TF U84 ( .A0(N312), .A1(DIVISION_HEAD[2]), .A2(N736), .B0(N311), .B1(
        N312), .Y(N313) );
  OAI2BB1X2TF U85 ( .A0N(N88), .A1N(C152_DATA4_11), .B0(N193), .Y(N936) );
  INVX2TF U86 ( .A(X_IN[5]), .Y(N60) );
  AND2X8TF U87 ( .A(N205), .B(ALU_START), .Y(N969) );
  CLKINVX4TF U88 ( .A(N969), .Y(N81) );
  INVX2TF U89 ( .A(X_IN[3]), .Y(N55) );
  AOI2BB1X4TF U90 ( .A0N(N961), .A1N(N960), .B0(N959), .Y(N1010) );
  OA21XLTF U91 ( .A0(SUM_AB[12]), .A1(N395), .B0(N73), .Y(N41) );
  INVX2TF U92 ( .A(N123), .Y(N46) );
  AOI22X1TF U93 ( .A0(N95), .A1(\INTADD_0_SUM[2] ), .B0(SUM_AB[3]), .B1(N85), 
        .Y(N423) );
  AOI22X1TF U94 ( .A0(N95), .A1(\INTADD_0_SUM[1] ), .B0(SUM_AB[2]), .B1(N85), 
        .Y(N413) );
  INVX2TF U95 ( .A(N1018), .Y(N49) );
  NOR2X1TF U96 ( .A(SUM_AB[8]), .B(N463), .Y(N478) );
  OR2X2TF U97 ( .A(N1010), .B(N82), .Y(N1011) );
  NOR2X1TF U98 ( .A(OPER_A[9]), .B(N900), .Y(N913) );
  OAI31X2TF U99 ( .A0(XTEMP[12]), .A1(N357), .A2(N511), .B0(N354), .Y(N355) );
  CLKINVX1TF U100 ( .A(SUM_AB[4]), .Y(N390) );
  AOI22X1TF U101 ( .A0(DIVISION_HEAD[1]), .A1(N72), .B0(ZTEMP[10]), .B1(N46), 
        .Y(N239) );
  OR2X2TF U102 ( .A(N348), .B(N599), .Y(N811) );
  INVX6TF U103 ( .A(DP_OP_333_124_4748_N57), .Y(N94) );
  OR2X2TF U104 ( .A(N142), .B(N228), .Y(N241) );
  CLKAND2X2TF U105 ( .A(ZTEMP[0]), .B(N244), .Y(POUT[0]) );
  AND2X6TF U106 ( .A(N178), .B(ALU_TYPE[1]), .Y(N205) );
  NAND2XLTF U107 ( .A(DIVISION_HEAD[4]), .B(N245), .Y(N207) );
  BUFX6TF U108 ( .A(X_IN[2]), .Y(N174) );
  CLKINVX1TF U109 ( .A(Y_IN[6]), .Y(N180) );
  AOI211X1TF U110 ( .A0(N56), .A1(N745), .B0(N441), .C0(N440), .Y(N442) );
  AOI211X1TF U111 ( .A0(Y_IN[7]), .A1(N745), .B0(N785), .C0(N784), .Y(N786) );
  AOI211X1TF U112 ( .A0(N61), .A1(N745), .B0(N459), .C0(N458), .Y(N460) );
  AOI22X1TF U113 ( .A0(N95), .A1(\INTADD_0_SUM[3] ), .B0(SUM_AB[4]), .B1(N85), 
        .Y(N432) );
  AOI22X1TF U114 ( .A0(N509), .A1(N466), .B0(SUM_AB[8]), .B1(N84), .Y(N468) );
  AOI22X1TF U115 ( .A0(N509), .A1(\INTADD_0_SUM[0] ), .B0(SUM_AB[1]), .B1(N85), 
        .Y(N403) );
  AOI22X1TF U116 ( .A0(N95), .A1(\INTADD_0_SUM[6] ), .B0(SUM_AB[7]), .B1(N85), 
        .Y(N462) );
  AOI22X1TF U117 ( .A0(N509), .A1(\INTADD_0_SUM[4] ), .B0(SUM_AB[5]), .B1(N84), 
        .Y(N439) );
  NAND2X1TF U118 ( .A(N500), .B(N499), .Y(N1013) );
  NOR2X1TF U119 ( .A(SUM_AB[10]), .B(N487), .Y(N500) );
  AOI21X1TF U120 ( .A0(SUM_AB[8]), .A1(N463), .B0(N478), .Y(N997) );
  NAND2X1TF U121 ( .A(N478), .B(N477), .Y(N487) );
  NOR2X4TF U122 ( .A(N920), .B(N912), .Y(N928) );
  NAND2X1TF U123 ( .A(N911), .B(N913), .Y(N930) );
  NAND2X1TF U124 ( .A(N454), .B(N453), .Y(N463) );
  NOR2X1TF U125 ( .A(SUM_AB[6]), .B(N444), .Y(N454) );
  NAND2X1TF U126 ( .A(N434), .B(N433), .Y(N444) );
  INVX4TF U127 ( .A(N767), .Y(N557) );
  NAND2X1TF U128 ( .A(N885), .B(N886), .Y(N900) );
  NOR2X1TF U129 ( .A(SUM_AB[4]), .B(N424), .Y(N434) );
  NAND2X1TF U130 ( .A(N416), .B(N415), .Y(N424) );
  NAND2X1TF U131 ( .A(N864), .B(N865), .Y(N879) );
  ADDHX2TF U132 ( .A(DP_OP_333_124_4748_N25), .B(DP_OP_333_124_4748_N9), .CO(
        DP_OP_333_124_4748_N8), .S(C152_DATA4_4) );
  OAI21X1TF U133 ( .A0(N379), .A1(N745), .B0(N381), .Y(N380) );
  NAND2X1TF U134 ( .A(N852), .B(N845), .Y(N855) );
  NOR3X1TF U135 ( .A(SUM_AB[0]), .B(SUM_AB[2]), .C(SUM_AB[1]), .Y(N416) );
  INVX1TF U136 ( .A(N405), .Y(N406) );
  AOI22X1TF U137 ( .A0(N174), .A1(N66), .B0(N56), .B1(N83), .Y(N783) );
  AOI22X1TF U138 ( .A0(Y_IN[9]), .A1(N800), .B0(N175), .B1(N66), .Y(N801) );
  AOI22X1TF U139 ( .A0(X_IN[12]), .A1(N83), .B0(X_IN[11]), .B1(N66), .Y(N437)
         );
  AOI22X1TF U140 ( .A0(DIVISION_HEAD[6]), .A1(N502), .B0(N176), .B1(N66), .Y(
        N399) );
  AOI32X1TF U141 ( .A0(N78), .A1(N45), .A2(N563), .B0(N617), .B1(N64), .Y(N544) );
  NAND3XLTF U142 ( .A(N78), .B(N822), .C(N821), .Y(N632) );
  OAI2BB2XLTF U143 ( .B0(N759), .B1(N802), .A0N(Y_IN[6]), .A1N(N800), .Y(N776)
         );
  OAI31XLTF U144 ( .A0(N75), .A1(N120), .A2(N631), .B0(N630), .Y(N636) );
  AOI22X1TF U145 ( .A0(XTEMP[10]), .A1(N99), .B0(N176), .B1(N800), .Y(N481) );
  NOR3X1TF U146 ( .A(OPER_A[2]), .B(OPER_A[1]), .C(OPER_A[0]), .Y(N838) );
  NOR2X1TF U147 ( .A(OPER_B[9]), .B(N899), .Y(N919) );
  OAI211XLTF U148 ( .A0(N81), .A1(N365), .B0(N971), .C0(N600), .Y(N367) );
  CLKINVX2TF U149 ( .A(OPER_A[0]), .Y(N829) );
  INVX1TF U150 ( .A(OPER_A[1]), .Y(N830) );
  INVX1TF U151 ( .A(OPER_A[11]), .Y(N927) );
  NAND2X1TF U152 ( .A(N883), .B(N139), .Y(N899) );
  OAI21X1TF U153 ( .A0(N126), .A1(N48), .B0(N231), .Y(OPER_A[2]) );
  OAI21X2TF U154 ( .A0(N119), .A1(N48), .B0(N230), .Y(OPER_A[1]) );
  OR2X2TF U155 ( .A(N387), .B(N766), .Y(N805) );
  OR2X2TF U156 ( .A(N387), .B(N761), .Y(N799) );
  AOI22X1TF U157 ( .A0(DIVISION_REMA[3]), .A1(N71), .B0(ZTEMP[3]), .B1(N142), 
        .Y(N232) );
  AOI22X1TF U158 ( .A0(DIVISION_HEAD[3]), .A1(N72), .B0(ZTEMP[12]), .B1(N46), 
        .Y(N242) );
  AOI22X1TF U159 ( .A0(DIVISION_REMA[4]), .A1(N72), .B0(ZTEMP[4]), .B1(N142), 
        .Y(N233) );
  AOI22X1TF U160 ( .A0(DIVISION_REMA[6]), .A1(N72), .B0(ZTEMP[6]), .B1(N142), 
        .Y(N235) );
  INVX2TF U161 ( .A(N745), .Y(N58) );
  AOI22X1TF U162 ( .A0(DIVISION_REMA[5]), .A1(N72), .B0(ZTEMP[5]), .B1(N142), 
        .Y(N234) );
  AOI22X1TF U163 ( .A0(DIVISION_REMA[1]), .A1(N71), .B0(ZTEMP[1]), .B1(N142), 
        .Y(N230) );
  NAND2X2TF U164 ( .A(N384), .B(N351), .Y(N734) );
  AOI22X1TF U165 ( .A0(DIVISION_REMA[0]), .A1(N71), .B0(ZTEMP[0]), .B1(N142), 
        .Y(N229) );
  AOI22X1TF U166 ( .A0(DIVISION_REMA[7]), .A1(N72), .B0(ZTEMP[7]), .B1(N142), 
        .Y(N236) );
  AOI22X1TF U167 ( .A0(DIVISION_REMA[8]), .A1(N72), .B0(ZTEMP[8]), .B1(N142), 
        .Y(N237) );
  AOI22X1TF U168 ( .A0(DIVISION_HEAD[0]), .A1(N72), .B0(ZTEMP[9]), .B1(N46), 
        .Y(N238) );
  AOI22X1TF U169 ( .A0(DIVISION_REMA[2]), .A1(N71), .B0(ZTEMP[2]), .B1(N142), 
        .Y(N231) );
  NOR2X1TF U170 ( .A(N858), .B(OPER_B[6]), .Y(N875) );
  INVX2TF U171 ( .A(N811), .Y(N76) );
  INVX8TF U172 ( .A(DP_OP_333_124_4748_N57), .Y(N185) );
  AND2X2TF U173 ( .A(N335), .B(N204), .Y(N944) );
  CLKINVX2TF U174 ( .A(N335), .Y(N953) );
  NAND2X2TF U175 ( .A(N353), .B(N306), .Y(N802) );
  AND2X2TF U176 ( .A(N351), .B(DP_OP_333_124_4748_N57), .Y(N745) );
  NAND2XLTF U177 ( .A(N204), .B(N948), .Y(N533) );
  AND2X2TF U178 ( .A(N123), .B(N228), .Y(N243) );
  NAND2X1TF U179 ( .A(N848), .B(N155), .Y(N854) );
  AND2X6TF U180 ( .A(ALU_START), .B(N244), .Y(N204) );
  OAI31X1TF U181 ( .A0(N965), .A1(N45), .A2(N970), .B0(N964), .Y(N966) );
  NAND2X1TF U182 ( .A(N156), .B(N365), .Y(N348) );
  AOI31X1TF U183 ( .A0(N157), .A1(N45), .A2(N963), .B0(N962), .Y(N964) );
  NOR2X1TF U184 ( .A(SIGN_Y), .B(N65), .Y(N896) );
  NAND2XLTF U185 ( .A(N605), .B(N822), .Y(N337) );
  NOR2X1TF U186 ( .A(OPER_B[3]), .B(N837), .Y(N848) );
  NAND2X1TF U187 ( .A(N124), .B(N305), .Y(N365) );
  AOI22X1TF U188 ( .A0(N64), .A1(DIVISION_HEAD[3]), .B0(XTEMP[12]), .B1(N45), 
        .Y(N342) );
  AND2X2TF U189 ( .A(N244), .B(N64), .Y(N225) );
  AND2X1TF U190 ( .A(ZTEMP[4]), .B(N244), .Y(POUT[4]) );
  AND2X2TF U191 ( .A(N65), .B(N244), .Y(N226) );
  OAI211X1TF U192 ( .A0(Y_IN[2]), .A1(N43), .B0(N310), .C0(N309), .Y(N311) );
  AND2X1TF U193 ( .A(ZTEMP[1]), .B(N244), .Y(POUT[1]) );
  INVX2TF U194 ( .A(N64), .Y(N65) );
  OR2X1TF U195 ( .A(N631), .B(N147), .Y(N369) );
  CLKINVX1TF U196 ( .A(N620), .Y(N622) );
  NAND2X1TF U197 ( .A(N834), .B(N154), .Y(N837) );
  INVX2TF U198 ( .A(Y_IN[7]), .Y(N173) );
  INVX8TF U199 ( .A(X_IN[0]), .Y(N747) );
  INVX2TF U200 ( .A(X_IN[11]), .Y(N177) );
  INVX2TF U201 ( .A(N501), .Y(N50) );
  INVX6TF U202 ( .A(Y_IN[1]), .Y(N307) );
  AOI21X2TF U203 ( .A0(N57), .A1(N42), .B0(N321), .Y(N323) );
  NOR3BX4TF U204 ( .AN(ALU_TYPE[0]), .B(ALU_TYPE[1]), .C(ALU_TYPE[2]), .Y(N244) );
  INVX2TF U205 ( .A(N226), .Y(N51) );
  INVX2TF U206 ( .A(N226), .Y(N52) );
  INVX2TF U207 ( .A(N225), .Y(N53) );
  INVX2TF U208 ( .A(N225), .Y(N54) );
  INVX2TF U209 ( .A(N55), .Y(N56) );
  INVX2TF U210 ( .A(N173), .Y(N57) );
  AOI32X4TF U211 ( .A0(N968), .A1(N967), .A2(N966), .B0(N78), .B1(N967), .Y(
        N1018) );
  INVX2TF U212 ( .A(N745), .Y(N59) );
  INVX2TF U213 ( .A(N60), .Y(N61) );
  INVX2TF U214 ( .A(N396), .Y(N62) );
  INVX2TF U215 ( .A(N396), .Y(N63) );
  INVX2TF U216 ( .A(N799), .Y(N66) );
  INVX2TF U217 ( .A(N799), .Y(N67) );
  INVX2TF U218 ( .A(N1011), .Y(N68) );
  INVX2TF U219 ( .A(N1011), .Y(N69) );
  INVX2TF U220 ( .A(N243), .Y(N70) );
  INVX2TF U221 ( .A(N241), .Y(N71) );
  INVX2TF U222 ( .A(N241), .Y(N72) );
  INVX2TF U223 ( .A(N944), .Y(N73) );
  INVX2TF U224 ( .A(N944), .Y(N75) );
  INVX2TF U225 ( .A(N811), .Y(N77) );
  INVX2TF U226 ( .A(N73), .Y(N78) );
  INVX2TF U227 ( .A(N47), .Y(N79) );
  INVX2TF U228 ( .A(N47), .Y(N80) );
  INVX2TF U229 ( .A(N969), .Y(N82) );
  INVX2TF U230 ( .A(N805), .Y(N83) );
  INVX2TF U231 ( .A(N41), .Y(N84) );
  INVX2TF U232 ( .A(N41), .Y(N85) );
  AOI22X1TF U233 ( .A0(N64), .A1(N141), .B0(POST_WORK), .B1(N65), .Y(N228) );
  NAND2X2TF U234 ( .A(N123), .B(N760), .Y(N455) );
  INVX2TF U235 ( .A(N177), .Y(N86) );
  CLKBUFX2TF U236 ( .A(Y_IN[5]), .Y(N172) );
  OAI22XLTF U237 ( .A0(N119), .A1(N734), .B0(N126), .B1(N455), .Y(N407) );
  OAI22XLTF U238 ( .A0(N42), .A1(N734), .B0(N130), .B1(N455), .Y(N430) );
  CLKBUFX2TF U239 ( .A(N227), .Y(N87) );
  NOR3BX1TF U240 ( .AN(ALU_TYPE[2]), .B(ALU_TYPE[0]), .C(ALU_TYPE[1]), .Y(N245) );
  CLKBUFX2TF U241 ( .A(N200), .Y(N88) );
  NAND2X1TF U242 ( .A(C152_DATA4_12), .B(N88), .Y(N202) );
  INVX2TF U243 ( .A(N898), .Y(N89) );
  NAND2X4TF U244 ( .A(N892), .B(N918), .Y(N934) );
  NOR2X6TF U245 ( .A(N203), .B(N75), .Y(N892) );
  CLKBUFX2TF U246 ( .A(DP_OP_333_124_4748_N43), .Y(N93) );
  OAI2BB2XLTF U247 ( .B0(OFFSET[0]), .B1(N185), .A0N(Y_IN[2]), .A1N(
        DP_OP_333_124_4748_N43), .Y(C2_Z_2) );
  AOI22XLTF U248 ( .A0(N172), .A1(N800), .B0(Y_IN[7]), .B1(N788), .Y(N752) );
  AOI22XLTF U249 ( .A0(DIVISION_HEAD[2]), .A1(N77), .B0(Y_IN[8]), .B1(N800), 
        .Y(N792) );
  AOI22XLTF U250 ( .A0(Y_IN[1]), .A1(N800), .B0(DIVISION_REMA[4]), .B1(N77), 
        .Y(N730) );
  AOI22XLTF U251 ( .A0(Y_IN[3]), .A1(N800), .B0(DIVISION_REMA[6]), .B1(N77), 
        .Y(N740) );
  NOR4XLTF U252 ( .A(N760), .B(N617), .C(N800), .D(N647), .Y(N248) );
  INVX2TF U253 ( .A(N511), .Y(N95) );
  AOI32X1TF U254 ( .A0(N509), .A1(DIVISION_HEAD[4]), .A2(N747), .B0(N472), 
        .B1(DIVISION_HEAD[4]), .Y(N393) );
  AOI21X2TF U255 ( .A0(N774), .A1(N373), .B0(N821), .Y(N509) );
  INVX2TF U256 ( .A(N967), .Y(N96) );
  AOI211X1TF U257 ( .A0(OPER_A[11]), .A1(N938), .B0(N937), .C0(N936), .Y(N939)
         );
  OAI2BB2XLTF U258 ( .B0(N872), .B1(N970), .A0N(C152_DATA4_6), .A1N(N88), .Y(
        N196) );
  NAND2X2TF U259 ( .A(SIGN_Y), .B(N963), .Y(N970) );
  NAND2X4TF U260 ( .A(N968), .B(N925), .Y(N906) );
  AOI21X2TF U261 ( .A0(N950), .A1(N965), .B0(N363), .Y(N968) );
  NOR3X2TF U262 ( .A(N121), .B(N122), .C(N952), .Y(N820) );
  NAND2X2TF U263 ( .A(N760), .B(N46), .Y(N558) );
  AOI22XLTF U264 ( .A0(DIVISION_HEAD[2]), .A1(N72), .B0(ZTEMP[11]), .B1(N46), 
        .Y(N240) );
  NOR4X2TF U265 ( .A(N647), .B(N945), .C(N367), .D(N366), .Y(N641) );
  CLKBUFX2TF U266 ( .A(N797), .Y(N98) );
  OAI21X1TF U267 ( .A0(SUM_AB[12]), .A1(N649), .B0(N73), .Y(N797) );
  CLKBUFX2TF U268 ( .A(N502), .Y(N99) );
  NOR3X1TF U269 ( .A(PRE_WORK), .B(N605), .C(N599), .Y(N502) );
  CMPR22X4TF U270 ( .A(DP_OP_333_124_4748_N24), .B(DP_OP_333_124_4748_N8), 
        .CO(DP_OP_333_124_4748_N7), .S(C152_DATA4_5) );
  XNOR2X1TF U271 ( .A(OPER_A[12]), .B(ADD_X_132_1_N2), .Y(N100) );
  CMPR32X2TF U272 ( .A(OPER_A[8]), .B(OPER_B[8]), .C(ADD_X_132_1_N6), .CO(
        ADD_X_132_1_N5), .S(SUM_AB[8]) );
  XNOR2X2TF U273 ( .A(N100), .B(OPER_B[12]), .Y(SUM_AB[12]) );
  ADDHX1TF U274 ( .A(OPER_B[0]), .B(OPER_A[0]), .CO(ADD_X_132_1_N13), .S(
        SUM_AB[0]) );
  AOI32X1TF U275 ( .A0(N273), .A1(N272), .A2(N309), .B0(N271), .B1(N272), .Y(
        N274) );
  OAI32X2TF U276 ( .A0(N270), .A1(N175), .A2(N307), .B0(X_IN[3]), .B1(N270), 
        .Y(N273) );
  OAI32X2TF U277 ( .A0(N250), .A1(N174), .A2(N307), .B0(X_IN[1]), .B1(N250), 
        .Y(N252) );
  NOR3BX4TF U278 ( .AN(N386), .B(N383), .C(N79), .Y(N514) );
  OR2X4TF U279 ( .A(N926), .B(N874), .Y(N189) );
  NAND2BX4TF U280 ( .AN(N819), .B(N856), .Y(N874) );
  OAI22X2TF U281 ( .A0(Y_IN[12]), .A1(N135), .B0(N330), .B1(N329), .Y(N331) );
  OAI22X4TF U282 ( .A0(N514), .A1(N359), .B0(N358), .B1(N44), .Y(N723) );
  AOI211X2TF U283 ( .A0(N494), .A1(N1012), .B0(N356), .C0(N355), .Y(N359) );
  OAI32X4TF U284 ( .A0(N284), .A1(X_IN[3]), .A2(N307), .B0(N174), .B1(N284), 
        .Y(N287) );
  AO22X4TF U285 ( .A0(N175), .A1(N736), .B0(X_IN[3]), .B1(N308), .Y(N284) );
  OAI32X4TF U286 ( .A0(N765), .A1(N764), .A2(X_IN[0]), .B0(N763), .B1(N765), 
        .Y(N768) );
  AOI2BB1X2TF U287 ( .A0N(X_IN[1]), .A1N(N762), .B0(N761), .Y(N765) );
  XOR2X4TF U288 ( .A(X_IN[12]), .B(N352), .Y(N357) );
  AOI222X4TF U289 ( .A0(XTEMP[11]), .A1(X_IN[11]), .B0(XTEMP[11]), .B1(N498), 
        .C0(X_IN[11]), .C1(N498), .Y(N352) );
  OAI21X1TF U290 ( .A0(N303), .A1(N383), .B0(N619), .Y(N304) );
  AOI32X1TF U291 ( .A0(N1017), .A1(N1014), .A2(N1013), .B0(N1012), .B1(N1014), 
        .Y(N1015) );
  NAND2X1TF U292 ( .A(N88), .B(C152_DATA4_9), .Y(N191) );
  NAND3X2TF U293 ( .A(N248), .B(N361), .C(N633), .Y(N619) );
  NOR2BX2TF U294 ( .AN(N543), .B(N384), .Y(N628) );
  AOI22X2TF U295 ( .A0(N342), .A1(N337), .B0(N943), .B1(N343), .Y(N918) );
  NOR2X2TF U296 ( .A(N332), .B(N954), .Y(N351) );
  NOR2X1TF U297 ( .A(ALU_TYPE[2]), .B(ALU_TYPE[0]), .Y(N178) );
  OAI21X1TF U298 ( .A0(N973), .A1(N906), .B0(N835), .Y(N871) );
  OAI22XLTF U299 ( .A0(N131), .A1(N734), .B0(N443), .B1(N59), .Y(N451) );
  NAND2X1TF U300 ( .A(PRE_WORK), .B(DP_OP_333_124_4748_N43), .Y(N387) );
  NOR2X1TF U301 ( .A(N124), .B(N627), .Y(N333) );
  OAI32X1TF U302 ( .A0(N648), .A1(N157), .A2(N946), .B0(N40), .B1(N649), .Y(
        N694) );
  OAI2BB2XLTF U303 ( .B0(N869), .B1(N920), .A0N(N203), .A1N(OPER_B[6]), .Y(
        N870) );
  NOR2BX1TF U304 ( .AN(N875), .B(OPER_B[7]), .Y(N883) );
  NAND2X1TF U305 ( .A(N565), .B(N384), .Y(N609) );
  INVX2TF U306 ( .A(N599), .Y(N566) );
  INVX2TF U307 ( .A(Y_IN[9]), .Y(N781) );
  AOI21X4TF U308 ( .A0(Y_IN[7]), .A1(N489), .B0(N260), .Y(N261) );
  CLKBUFX2TF U309 ( .A(X_IN[7]), .Y(N176) );
  OAI21X1TF U310 ( .A0(N42), .A1(N48), .B0(N232), .Y(OPER_A[3]) );
  NAND2X1TF U311 ( .A(N122), .B(N147), .Y(N604) );
  NAND2X1TF U312 ( .A(N134), .B(N149), .Y(N332) );
  AOI211X2TF U313 ( .A0(N570), .A1(N78), .B0(N594), .C0(N569), .Y(N596) );
  NAND2X1TF U314 ( .A(N892), .B(N916), .Y(N941) );
  NAND3X2TF U315 ( .A(N202), .B(N346), .C(N201), .Y(N724) );
  OAI2BB1X1TF U316 ( .A0N(DIVISION_HEAD[10]), .A1N(N472), .B0(N452), .Y(N713)
         );
  OAI22X1TF U317 ( .A0(N75), .A1(N1017), .B0(N503), .B1(N59), .Y(N356) );
  CLKINVX6TF U318 ( .A(N892), .Y(N920) );
  OAI21X1TF U319 ( .A0(Y_IN[11]), .A1(N127), .B0(N322), .Y(N324) );
  NAND2X1TF U320 ( .A(N121), .B(N120), .Y(N603) );
  NAND3X1TF U321 ( .A(N960), .B(N82), .C(N599), .Y(N646) );
  INVX12TF U322 ( .A(Y_IN[3]), .Y(N729) );
  NAND2X6TF U323 ( .A(Y_IN[1]), .B(Y_IN[0]), .Y(N308) );
  INVX2TF U324 ( .A(X_IN[8]), .Y(N489) );
  AND2X8TF U325 ( .A(N204), .B(PRE_WORK), .Y(DP_OP_333_124_4748_N57) );
  AOI32X1TF U326 ( .A0(N565), .A1(N77), .A2(N161), .B0(N958), .B1(N76), .Y(
        N567) );
  NOR3X1TF U327 ( .A(N605), .B(N604), .C(N774), .Y(N606) );
  AOI222X2TF U328 ( .A0(DIVISION_HEAD[1]), .A1(DIVISION_HEAD[0]), .B0(
        DIVISION_HEAD[1]), .B1(N308), .C0(DIVISION_HEAD[0]), .C1(N307), .Y(
        N310) );
  NAND2X1TF U329 ( .A(N134), .B(STEP[3]), .Y(N631) );
  NAND2X1TF U330 ( .A(N121), .B(N122), .Y(N954) );
  NOR2X1TF U331 ( .A(N156), .B(N599), .Y(N353) );
  NAND2X2TF U332 ( .A(ALU_START), .B(N245), .Y(N599) );
  INVX2TF U333 ( .A(Y_IN[8]), .Y(N759) );
  INVX2TF U334 ( .A(Y_IN[10]), .Y(N547) );
  NOR2X2TF U335 ( .A(N348), .B(N81), .Y(N384) );
  OAI22X1TF U336 ( .A0(DIVISION_HEAD[12]), .A1(N144), .B0(XTEMP[12]), .B1(N40), 
        .Y(N537) );
  NAND4BX1TF U337 ( .AN(N824), .B(N827), .C(N195), .D(N194), .Y(N681) );
  AOI222X4TF U338 ( .A0(N488), .A1(N136), .B0(N488), .B1(N503), .C0(N136), 
        .C1(N503), .Y(N498) );
  NOR2X1TF U339 ( .A(OPER_B[5]), .B(N854), .Y(N862) );
  INVX2TF U340 ( .A(N1014), .Y(N1009) );
  AOI2BB1X1TF U341 ( .A0N(N607), .A1N(N336), .B0(N960), .Y(N179) );
  AOI2BB1X4TF U342 ( .A0N(DIVISION_HEAD[6]), .A1N(N320), .B0(Y_IN[6]), .Y(N318) );
  AOI2BB1X4TF U343 ( .A0N(DIVISION_HEAD[4]), .A1N(N316), .B0(Y_IN[4]), .Y(N314) );
  NOR2X1TF U344 ( .A(N172), .B(N119), .Y(N315) );
  NOR2X4TF U345 ( .A(Y_IN[3]), .B(N40), .Y(N312) );
  NOR2X2TF U346 ( .A(N760), .B(N170), .Y(N758) );
  NOR2X2TF U347 ( .A(\RSHT_BITS[3] ), .B(N591), .Y(N605) );
  AOI211X2TF U348 ( .A0(X_IN[10]), .A1(N759), .B0(N294), .C0(N293), .Y(N297)
         );
  AOI21X2TF U349 ( .A0(Y_IN[7]), .A1(N501), .B0(N292), .Y(N293) );
  AOI211X2TF U350 ( .A0(X_IN[8]), .A1(N291), .B0(N290), .C0(N289), .Y(N292) );
  AOI32X4TF U351 ( .A0(N287), .A1(N286), .A2(N309), .B0(N285), .B1(N286), .Y(
        N288) );
  OA21X4TF U352 ( .A0(N759), .A1(N86), .B0(N279), .Y(N281) );
  AOI21X2TF U353 ( .A0(Y_IN[7]), .A1(N503), .B0(N278), .Y(N279) );
  AOI211X2TF U354 ( .A0(X_IN[9]), .A1(N277), .B0(N276), .C0(N275), .Y(N278) );
  AO22X2TF U355 ( .A0(X_IN[5]), .A1(N736), .B0(N175), .B1(N308), .Y(N270) );
  AOI21X4TF U356 ( .A0(N172), .A1(N464), .B0(N256), .Y(N259) );
  OAI211X4TF U357 ( .A0(Y_IN[3]), .A1(N443), .B0(N249), .C0(N309), .Y(N250) );
  INVX6TF U358 ( .A(Y_IN[2]), .Y(N736) );
  INVX2TF U359 ( .A(X_IN[10]), .Y(N503) );
  OAI21X1TF U360 ( .A0(N131), .A1(N48), .B0(N234), .Y(OPER_A[5]) );
  NOR2X2TF U361 ( .A(N332), .B(N604), .Y(N958) );
  AOI211X1TF U362 ( .A0(N204), .A1(N607), .B0(N947), .C0(N606), .Y(N610) );
  NOR2X1TF U363 ( .A(N604), .B(N952), .Y(N564) );
  NAND2X1TF U364 ( .A(STEP[2]), .B(N149), .Y(N952) );
  INVX2TF U365 ( .A(N958), .Y(N965) );
  NAND2X1TF U366 ( .A(N896), .B(N74), .Y(N956) );
  NAND2X1TF U367 ( .A(N333), .B(N156), .Y(N338) );
  AOI21X4TF U368 ( .A0(Y_IN[3]), .A1(N40), .B0(N313), .Y(N316) );
  AOI31X1TF U369 ( .A0(N78), .A1(N64), .A2(N563), .B0(N350), .Y(N386) );
  NAND2X1TF U370 ( .A(N565), .B(DP_OP_333_124_4748_N57), .Y(N395) );
  NOR2X2TF U371 ( .A(N332), .B(N603), .Y(N565) );
  NAND3X1TF U372 ( .A(N92), .B(N91), .C(N90), .Y(N591) );
  INVX2TF U373 ( .A(N58), .Y(N800) );
  INVX2TF U374 ( .A(N204), .Y(N960) );
  AOI2BB1X2TF U375 ( .A0N(N291), .A1N(X_IN[8]), .B0(Y_IN[6]), .Y(N289) );
  NAND2X2TF U376 ( .A(X_IN[5]), .B(N729), .Y(N286) );
  NAND2X1TF U377 ( .A(MODE_TYPE[0]), .B(N306), .Y(N761) );
  NOR4X2TF U378 ( .A(Y_IN[12]), .B(Y_IN[11]), .C(Y_IN[10]), .D(N282), .Y(N283)
         );
  AOI211X2TF U379 ( .A0(N86), .A1(N759), .B0(N281), .C0(N280), .Y(N282) );
  AOI2BB1X2TF U380 ( .A0N(N277), .A1N(N50), .B0(Y_IN[6]), .Y(N275) );
  AOI211X2TF U381 ( .A0(X_IN[9]), .A1(N759), .B0(N262), .C0(N261), .Y(N266) );
  AOI211X2TF U382 ( .A0(N259), .A1(N176), .B0(N258), .C0(N257), .Y(N260) );
  AOI2BB1X2TF U383 ( .A0N(N176), .A1N(N259), .B0(Y_IN[6]), .Y(N257) );
  AOI211X2TF U384 ( .A0(N255), .A1(N61), .B0(N254), .C0(N253), .Y(N256) );
  AOI2BB1X2TF U385 ( .A0N(N61), .A1N(N255), .B0(Y_IN[4]), .Y(N253) );
  AOI211X4TF U386 ( .A0(Y_IN[3]), .A1(N443), .B0(N252), .C0(N251), .Y(N255) );
  INVX2TF U387 ( .A(N364), .Y(N760) );
  NAND2X1TF U388 ( .A(N384), .B(N958), .Y(N364) );
  AOI222X4TF U389 ( .A0(XTEMP[9]), .A1(X_IN[9]), .B0(XTEMP[9]), .B1(N479), 
        .C0(X_IN[9]), .C1(N479), .Y(N488) );
  AOI222X4TF U390 ( .A0(N135), .A1(N489), .B0(N135), .B1(N465), .C0(N489), 
        .C1(N465), .Y(N479) );
  NAND2X1TF U391 ( .A(N948), .B(DP_OP_333_124_4748_N57), .Y(N634) );
  INVX12TF U392 ( .A(N925), .Y(N203) );
  NAND3X1TF U393 ( .A(STEP[2]), .B(STEP[3]), .C(N642), .Y(N943) );
  AOI211X2TF U394 ( .A0(DIVISION_HEAD[8]), .A1(N759), .B0(N323), .C0(N324), 
        .Y(N330) );
  AOI211X2TF U395 ( .A0(N320), .A1(DIVISION_HEAD[6]), .B0(N319), .C0(N318), 
        .Y(N321) );
  AOI21X4TF U396 ( .A0(N172), .A1(N119), .B0(N317), .Y(N320) );
  AOI211X2TF U397 ( .A0(N316), .A1(DIVISION_HEAD[4]), .B0(N315), .C0(N314), 
        .Y(N317) );
  NOR3X1TF U398 ( .A(N771), .B(N79), .C(N556), .Y(N779) );
  NOR2X1TF U399 ( .A(N954), .B(N631), .Y(N563) );
  OA22X4TF U400 ( .A0(N766), .A1(N557), .B0(N761), .B1(N762), .Y(N302) );
  NAND2X1TF U401 ( .A(N958), .B(DP_OP_333_124_4748_N57), .Y(N649) );
  AO22X1TF U402 ( .A0(N372), .A1(XTEMP[12]), .B0(N360), .B1(N963), .Y(N722) );
  NAND2X1TF U403 ( .A(N642), .B(N77), .Y(N614) );
  AOI32X1TF U404 ( .A0(N965), .A1(N361), .A2(N956), .B0(N971), .B1(N361), .Y(
        N362) );
  INVX2TF U405 ( .A(N509), .Y(N511) );
  OAI2BB2XLTF U406 ( .B0(N45), .B1(N970), .A0N(N970), .A1N(N45), .Y(N972) );
  NAND2X1TF U407 ( .A(N82), .B(N94), .Y(N186) );
  OR2X8TF U408 ( .A(N959), .B(N179), .Y(N925) );
  OAI21X4TF U409 ( .A0(N949), .A1(N609), .B0(N646), .Y(N959) );
  OAI21X4TF U410 ( .A0(DIVISION_HEAD[12]), .A1(N548), .B0(N331), .Y(N949) );
  NAND2X6TF U411 ( .A(N546), .B(N386), .Y(N461) );
  OAI211X1TF U412 ( .A0(N958), .A1(N348), .B0(N566), .C0(N600), .Y(N349) );
  INVX2TF U413 ( .A(N76), .Y(N774) );
  NOR2BX4TF U414 ( .AN(N546), .B(N556), .Y(N812) );
  NAND2X1TF U415 ( .A(N351), .B(N76), .Y(N543) );
  AOI31X4TF U416 ( .A0(N122), .A1(N385), .A2(N384), .B0(N383), .Y(N546) );
  AOI21X4TF U417 ( .A0(N764), .A1(N302), .B0(N387), .Y(N383) );
  AOI211X4TF U418 ( .A0(Y_IN[11]), .A1(N298), .B0(Y_IN[12]), .C0(N269), .Y(
        N764) );
  OAI21X1TF U419 ( .A0(N156), .A1(N647), .B0(N646), .Y(N695) );
  AOI22X1TF U420 ( .A0(N542), .A1(N64), .B0(N541), .B1(N540), .Y(N707) );
  INVX2TF U421 ( .A(N542), .Y(N540) );
  OAI31X1TF U422 ( .A0(N539), .A1(N538), .A2(N537), .B0(N536), .Y(N541) );
  AOI211X1TF U423 ( .A0(N535), .A1(XTEMP[12]), .B0(N534), .C0(N533), .Y(N536)
         );
  OAI31X1TF U424 ( .A0(DIVISION_HEAD[1]), .A1(N532), .A2(N136), .B0(N531), .Y(
        N535) );
  AOI22X1TF U425 ( .A0(N530), .A1(N529), .B0(XTEMP[11]), .B1(N43), .Y(N531) );
  OAI22X1TF U426 ( .A0(DIVISION_HEAD[0]), .A1(N39), .B0(DIVISION_REMA[8]), 
        .B1(N135), .Y(N529) );
  INVX2TF U427 ( .A(N538), .Y(N530) );
  NOR2X1TF U428 ( .A(XTEMP[11]), .B(N43), .Y(N532) );
  OAI21X1TF U429 ( .A0(XTEMP[11]), .A1(N43), .B0(N528), .Y(N538) );
  AOI22X1TF U430 ( .A0(DIVISION_HEAD[0]), .A1(N39), .B0(DIVISION_HEAD[1]), 
        .B1(N136), .Y(N528) );
  AOI21X1TF U431 ( .A0(DIVISION_HEAD[11]), .A1(N146), .B0(N527), .Y(N539) );
  AOI211X1TF U432 ( .A0(DIVISION_REMA[6]), .A1(N132), .B0(N526), .C0(N525), 
        .Y(N527) );
  NOR2X1TF U433 ( .A(DIVISION_HEAD[11]), .B(N146), .Y(N525) );
  AOI21X1TF U434 ( .A0(DIVISION_HEAD[9]), .A1(N145), .B0(N523), .Y(N524) );
  AOI211X1TF U435 ( .A0(DIVISION_REMA[4]), .A1(N130), .B0(N522), .C0(N521), 
        .Y(N523) );
  NOR2X1TF U436 ( .A(DIVISION_HEAD[9]), .B(N145), .Y(N521) );
  AOI21X1TF U437 ( .A0(DIVISION_HEAD[7]), .A1(N143), .B0(N519), .Y(N520) );
  AOI211X1TF U438 ( .A0(N518), .A1(DIVISION_REMA[2]), .B0(N517), .C0(N516), 
        .Y(N519) );
  NOR2X1TF U439 ( .A(DIVISION_HEAD[7]), .B(N143), .Y(N517) );
  OAI21X1TF U440 ( .A0(DIVISION_HEAD[5]), .A1(N158), .B0(N515), .Y(N518) );
  OAI211X1TF U441 ( .A0(DIVISION_REMA[1]), .A1(N119), .B0(DIVISION_REMA[0]), 
        .C0(N125), .Y(N515) );
  AOI22X1TF U442 ( .A0(N596), .A1(N92), .B0(N580), .B1(N579), .Y(N703) );
  AOI211X1TF U443 ( .A0(N594), .A1(N137), .B0(N578), .C0(N788), .Y(N580) );
  AOI21X1TF U444 ( .A0(N577), .A1(N774), .B0(N159), .Y(N578) );
  OAI21X1TF U445 ( .A0(N381), .A1(N141), .B0(N380), .Y(N720) );
  OAI22X1TF U446 ( .A0(N75), .A1(N378), .B0(N761), .B1(N639), .Y(N379) );
  AOI21X1TF U447 ( .A0(N820), .A1(N375), .B0(N374), .Y(N377) );
  OAI211X1TF U448 ( .A0(N373), .A1(N821), .B0(N611), .C0(N639), .Y(N374) );
  OAI21X1TF U449 ( .A0(N135), .A1(N227), .B0(N224), .Y(FOUT[8]) );
  AOI21X1TF U450 ( .A0(N205), .A1(DIVISION_REMA[8]), .B0(N223), .Y(N224) );
  OAI22X1TF U451 ( .A0(N150), .A1(N52), .B0(N136), .B1(N53), .Y(N223) );
  AND2X2TF U452 ( .A(ZTEMP[8]), .B(N97), .Y(POUT[8]) );
  OAI21X1TF U453 ( .A0(N42), .A1(N87), .B0(N214), .Y(FOUT[3]) );
  AOI21X1TF U454 ( .A0(N205), .A1(DIVISION_REMA[3]), .B0(N213), .Y(N214) );
  OAI22X1TF U455 ( .A0(N131), .A1(N54), .B0(N145), .B1(N52), .Y(N213) );
  AND2X2TF U456 ( .A(ZTEMP[3]), .B(N97), .Y(POUT[3]) );
  AOI22X1TF U457 ( .A0(N203), .A1(OPER_B[8]), .B0(N892), .B1(N891), .Y(N198)
         );
  OAI21X1TF U458 ( .A0(N890), .A1(N139), .B0(N889), .Y(N891) );
  AOI211X1TF U459 ( .A0(N916), .A1(OPER_B[9]), .B0(N888), .C0(N887), .Y(N889)
         );
  OAI32X1TF U460 ( .A0(OPER_A[8]), .A1(N886), .A2(N912), .B0(N885), .B1(N884), 
        .Y(N887) );
  AOI21X1TF U461 ( .A0(N909), .A1(N886), .B0(N908), .Y(N884) );
  NOR3X1TF U462 ( .A(N907), .B(OPER_B[8]), .C(N883), .Y(N888) );
  AOI21X1TF U463 ( .A0(N883), .A1(N918), .B0(N917), .Y(N890) );
  OAI21X1TF U464 ( .A0(N130), .A1(N227), .B0(N216), .Y(FOUT[4]) );
  AOI21X1TF U465 ( .A0(N205), .A1(DIVISION_REMA[4]), .B0(N215), .Y(N216) );
  OAI22X1TF U466 ( .A0(N132), .A1(N53), .B0(N152), .B1(N51), .Y(N215) );
  OAI21X1TF U467 ( .A0(N127), .A1(N227), .B0(N222), .Y(FOUT[7]) );
  AOI21X1TF U468 ( .A0(N205), .A1(DIVISION_REMA[7]), .B0(N221), .Y(N222) );
  OAI22X1TF U469 ( .A0(N148), .A1(N52), .B0(N39), .B1(N53), .Y(N221) );
  AND2X2TF U470 ( .A(ZTEMP[7]), .B(N97), .Y(POUT[7]) );
  OAI21X1TF U471 ( .A0(N596), .A1(N585), .B0(N584), .Y(N702) );
  AOI31X1TF U472 ( .A0(N583), .A1(N588), .A2(N590), .B0(N582), .Y(N585) );
  OAI22X1TF U473 ( .A0(N128), .A1(N581), .B0(N592), .B1(N588), .Y(N582) );
  AOI211X1TF U474 ( .A0(N203), .A1(OPER_B[10]), .B0(N923), .C0(N924), .Y(N199)
         );
  AOI21X1TF U475 ( .A0(N973), .A1(N970), .B0(N906), .Y(N924) );
  AOI21X1TF U476 ( .A0(N922), .A1(N921), .B0(N920), .Y(N923) );
  AOI32X1TF U477 ( .A0(N919), .A1(OPER_B[10]), .A2(N918), .B0(N917), .B1(
        OPER_B[10]), .Y(N921) );
  AOI211X1TF U478 ( .A0(N916), .A1(OPER_B[11]), .B0(N915), .C0(N914), .Y(N922)
         );
  OAI32X1TF U479 ( .A0(OPER_A[10]), .A1(N913), .A2(N912), .B0(N911), .B1(N910), 
        .Y(N914) );
  AOI21X1TF U480 ( .A0(N909), .A1(N913), .B0(N908), .Y(N910) );
  NOR3X1TF U481 ( .A(N907), .B(OPER_B[10]), .C(N919), .Y(N915) );
  OAI22X1TF U482 ( .A0(N90), .A1(N597), .B0(N596), .B1(N595), .Y(N701) );
  AOI21X1TF U483 ( .A0(\INDEX[2] ), .A1(N594), .B0(N593), .Y(N595) );
  OAI22X1TF U484 ( .A0(N592), .A1(N591), .B0(N590), .B1(N589), .Y(N593) );
  INVX2TF U485 ( .A(N587), .Y(N592) );
  AOI21X1TF U486 ( .A0(N588), .A1(N587), .B0(N586), .Y(N597) );
  OAI22X1TF U487 ( .A0(N596), .A1(N576), .B0(N575), .B1(N169), .Y(N704) );
  AOI21X1TF U488 ( .A0(N591), .A1(N587), .B0(N586), .Y(N575) );
  OAI21X1TF U489 ( .A0(N90), .A1(N590), .B0(N583), .Y(N589) );
  INVX2TF U490 ( .A(N614), .Y(N583) );
  INVX2TF U491 ( .A(N596), .Y(N579) );
  OAI31X1TF U492 ( .A0(N605), .A1(N604), .A2(N774), .B0(N577), .Y(N587) );
  OAI32X1TF U493 ( .A0(N574), .A1(N822), .A2(N573), .B0(N78), .B1(N574), .Y(
        N577) );
  INVX2TF U494 ( .A(N572), .Y(N574) );
  AOI21X1TF U495 ( .A0(N594), .A1(N166), .B0(N571), .Y(N576) );
  AOI31X1TF U496 ( .A0(N78), .A1(N822), .A2(N821), .B0(N946), .Y(N568) );
  INVX2TF U497 ( .A(N581), .Y(N594) );
  OAI31X1TF U498 ( .A0(N564), .A1(N565), .A2(N563), .B0(N78), .Y(N581) );
  OAI21X1TF U499 ( .A0(N129), .A1(N619), .B0(N304), .Y(N726) );
  AOI32X1TF U500 ( .A0(N628), .A1(N634), .A2(N376), .B0(N137), .B1(N634), .Y(
        N303) );
  AND2X2TF U501 ( .A(ZTEMP[10]), .B(N97), .Y(POUT[10]) );
  AND2X2TF U502 ( .A(ZTEMP[9]), .B(N97), .Y(POUT[9]) );
  OAI211X1TF U503 ( .A0(N1018), .A1(N1017), .B0(N1016), .C0(N1015), .Y(N657)
         );
  AOI22X1TF U504 ( .A0(DIVISION_HEAD[12]), .A1(N69), .B0(ZTEMP[12]), .B1(N1010), .Y(N1016) );
  OAI21X1TF U505 ( .A0(N132), .A1(N227), .B0(N220), .Y(FOUT[6]) );
  AOI21X1TF U506 ( .A0(N205), .A1(DIVISION_REMA[6]), .B0(N219), .Y(N220) );
  OAI22X1TF U507 ( .A0(N135), .A1(N54), .B0(N144), .B1(N51), .Y(N219) );
  AND2X2TF U508 ( .A(ZTEMP[6]), .B(N97), .Y(POUT[6]) );
  OAI21X1TF U509 ( .A0(N131), .A1(N227), .B0(N218), .Y(FOUT[5]) );
  AOI21X1TF U510 ( .A0(N205), .A1(DIVISION_REMA[5]), .B0(N217), .Y(N218) );
  OAI22X1TF U511 ( .A0(N127), .A1(N54), .B0(N146), .B1(N51), .Y(N217) );
  AND2X2TF U512 ( .A(ZTEMP[5]), .B(N97), .Y(POUT[5]) );
  NOR2X1TF U513 ( .A(N87), .B(N133), .Y(FOUT[11]) );
  AND2X2TF U514 ( .A(ZTEMP[11]), .B(N97), .Y(POUT[11]) );
  NOR2X1TF U515 ( .A(N87), .B(N44), .Y(FOUT[12]) );
  AND2X2TF U516 ( .A(ZTEMP[12]), .B(N97), .Y(POUT[12]) );
  INVX2TF U517 ( .A(N895), .Y(N872) );
  AOI211X1TF U518 ( .A0(OPER_B[6]), .A1(N868), .B0(N867), .C0(N866), .Y(N869)
         );
  OAI32X1TF U519 ( .A0(OPER_A[6]), .A1(N865), .A2(N912), .B0(N864), .B1(N863), 
        .Y(N866) );
  AOI21X1TF U520 ( .A0(N909), .A1(N865), .B0(N908), .Y(N863) );
  INVX2TF U521 ( .A(N912), .Y(N909) );
  OAI31X1TF U522 ( .A0(N907), .A1(OPER_B[6]), .A2(N862), .B0(N861), .Y(N867)
         );
  AOI21X1TF U523 ( .A0(OPER_B[7]), .A1(N860), .B0(N859), .Y(N861) );
  OAI21X1TF U524 ( .A0(N907), .A1(N858), .B0(N857), .Y(N868) );
  OAI21X1TF U525 ( .A0(N126), .A1(N227), .B0(N212), .Y(FOUT[2]) );
  AOI21X1TF U526 ( .A0(N205), .A1(DIVISION_REMA[2]), .B0(N211), .Y(N212) );
  OAI22X1TF U527 ( .A0(N130), .A1(N53), .B0(N151), .B1(N51), .Y(N211) );
  AND2X2TF U528 ( .A(ZTEMP[2]), .B(N97), .Y(POUT[2]) );
  OAI22X1TF U529 ( .A0(N514), .A1(N486), .B0(N485), .B1(N39), .Y(N710) );
  AOI211X1TF U530 ( .A0(SUM_AB[9]), .A1(N85), .B0(N483), .C0(N482), .Y(N486)
         );
  OAI211X1TF U531 ( .A0(N1002), .A1(N507), .B0(N481), .C0(N480), .Y(N482) );
  OAI22X1TF U532 ( .A0(N135), .A1(N47), .B0(N489), .B1(N608), .Y(N483) );
  AOI22X1TF U533 ( .A0(OPER_B[9]), .A1(N902), .B0(OPER_A[9]), .B1(N901), .Y(
        N903) );
  OAI21X1TF U534 ( .A0(N931), .A1(N900), .B0(N929), .Y(N901) );
  OAI21X1TF U535 ( .A0(N934), .A1(N899), .B0(N932), .Y(N902) );
  AOI31X1TF U536 ( .A0(N898), .A1(N168), .A2(N899), .B0(N897), .Y(N904) );
  OAI211X1TF U537 ( .A0(N140), .A1(N941), .B0(N191), .C0(N190), .Y(N897) );
  AOI22X1TF U538 ( .A0(SIGN_Y), .A1(N895), .B0(N894), .B1(N900), .Y(N905) );
  NOR2X1TF U539 ( .A(N931), .B(OPER_A[9]), .Y(N894) );
  OAI22X1TF U540 ( .A0(N514), .A1(N497), .B0(N496), .B1(N136), .Y(N709) );
  AOI21X1TF U541 ( .A0(N494), .A1(N1003), .B0(N493), .Y(N497) );
  OAI211X1TF U542 ( .A0(N501), .A1(N608), .B0(N492), .C0(N491), .Y(N493) );
  OAI22X1TF U543 ( .A0(N39), .A1(N734), .B0(N489), .B1(N58), .Y(N490) );
  AOI22X1TF U544 ( .A0(XTEMP[11]), .A1(N99), .B0(SUM_AB[10]), .B1(N84), .Y(
        N492) );
  OAI21X1TF U545 ( .A0(N758), .A1(N161), .B0(N562), .Y(N705) );
  OAI22X1TF U546 ( .A0(N561), .A1(N560), .B0(N760), .B1(N777), .Y(N562) );
  AOI22X1TF U547 ( .A0(Y_IN[0]), .A1(N788), .B0(DIVISION_REMA[1]), .B1(N77), 
        .Y(N559) );
  AOI21X1TF U548 ( .A0(N75), .A1(N649), .B0(N974), .Y(N561) );
  OAI21X1TF U549 ( .A0(N119), .A1(N227), .B0(N210), .Y(FOUT[1]) );
  AOI21X1TF U550 ( .A0(N205), .A1(DIVISION_REMA[1]), .B0(N209), .Y(N210) );
  OAI22X1TF U551 ( .A0(N42), .A1(N53), .B0(N143), .B1(N51), .Y(N209) );
  INVX2TF U552 ( .A(N245), .Y(N227) );
  OAI211X1TF U553 ( .A0(SIGN_Y), .A1(N963), .B0(N206), .C0(N970), .Y(N893) );
  OAI21X1TF U554 ( .A0(N128), .A1(N619), .B0(N618), .Y(N699) );
  AOI31X1TF U555 ( .A0(N617), .A1(N620), .A2(N616), .B0(N615), .Y(N618) );
  OAI32X1TF U556 ( .A0(N628), .A1(N629), .A2(N620), .B0(N616), .B1(N628), .Y(
        N615) );
  OAI22X1TF U557 ( .A0(N170), .A1(N739), .B0(N758), .B1(N151), .Y(N690) );
  AOI211X1TF U558 ( .A0(SUM_AB[4]), .A1(N98), .B0(N738), .C0(N737), .Y(N739)
         );
  OAI211X1TF U559 ( .A0(N736), .A1(N59), .B0(N754), .C0(N735), .Y(N737) );
  AOI22X1TF U560 ( .A0(DIVISION_REMA[5]), .A1(N77), .B0(N794), .B1(N985), .Y(
        N735) );
  OAI22X1TF U561 ( .A0(N182), .A1(N802), .B0(N143), .B1(N734), .Y(N738) );
  OAI22X1TF U562 ( .A0(N170), .A1(N728), .B0(N758), .B1(N153), .Y(N692) );
  AOI211X1TF U563 ( .A0(SUM_AB[2]), .A1(N98), .B0(N727), .C0(N656), .Y(N728)
         );
  OAI211X1TF U564 ( .A0(N655), .A1(N59), .B0(N754), .C0(N654), .Y(N656) );
  AOI22X1TF U565 ( .A0(DIVISION_REMA[3]), .A1(N77), .B0(N794), .B1(N979), .Y(
        N654) );
  OAI22X1TF U566 ( .A0(N736), .A1(N802), .B0(N158), .B1(N734), .Y(N727) );
  OAI22X1TF U567 ( .A0(N170), .A1(N653), .B0(N758), .B1(N158), .Y(N693) );
  AOI21X1TF U568 ( .A0(SUM_AB[1]), .A1(N98), .B0(N652), .Y(N653) );
  AOI22X1TF U569 ( .A0(DIVISION_REMA[0]), .A1(N80), .B0(N794), .B1(N976), .Y(
        N650) );
  AOI22X1TF U570 ( .A0(Y_IN[1]), .A1(N788), .B0(DIVISION_REMA[2]), .B1(N77), 
        .Y(N651) );
  OAI22X1TF U571 ( .A0(N170), .A1(N750), .B0(N758), .B1(N152), .Y(N688) );
  AOI211X1TF U572 ( .A0(N991), .A1(N794), .B0(N749), .C0(N748), .Y(N750) );
  OAI211X1TF U573 ( .A0(N747), .A1(N805), .B0(N754), .C0(N746), .Y(N748) );
  AOI22X1TF U574 ( .A0(DIVISION_REMA[7]), .A1(N76), .B0(SUM_AB[6]), .B1(N797), 
        .Y(N746) );
  OAI21X1TF U575 ( .A0(N182), .A1(N59), .B0(N744), .Y(N749) );
  AOI22X1TF U576 ( .A0(Y_IN[6]), .A1(N788), .B0(DIVISION_REMA[5]), .B1(N80), 
        .Y(N744) );
  OAI211X1TF U577 ( .A0(N167), .A1(N941), .B0(N940), .C0(N939), .Y(N671) );
  AOI21X1TF U578 ( .A0(N962), .A1(N206), .B0(N192), .Y(N193) );
  NOR3X1TF U579 ( .A(N934), .B(OPER_B[11]), .C(N935), .Y(N192) );
  INVX2TF U580 ( .A(N933), .Y(N935) );
  OAI32X1TF U581 ( .A0(N165), .A1(N933), .A2(N89), .B0(N932), .B1(N165), .Y(
        N937) );
  OAI21X1TF U582 ( .A0(N931), .A1(N930), .B0(N929), .Y(N938) );
  AOI31X1TF U583 ( .A0(N928), .A1(N927), .A2(N930), .B0(N926), .Y(N940) );
  AOI22X1TF U584 ( .A0(SUM_AB[10]), .A1(N171), .B0(N1003), .B1(N1014), .Y(
        N1004) );
  AOI22X1TF U585 ( .A0(DIVISION_HEAD[10]), .A1(N69), .B0(ZTEMP[10]), .B1(N96), 
        .Y(N1005) );
  AOI22X1TF U586 ( .A0(SUM_AB[8]), .A1(N171), .B0(N997), .B1(N1014), .Y(N998)
         );
  AOI22X1TF U587 ( .A0(DIVISION_HEAD[8]), .A1(N69), .B0(ZTEMP[8]), .B1(N96), 
        .Y(N999) );
  AOI22X1TF U588 ( .A0(SUM_AB[4]), .A1(N171), .B0(N985), .B1(N1014), .Y(N986)
         );
  AOI22X1TF U589 ( .A0(DIVISION_HEAD[4]), .A1(N69), .B0(ZTEMP[4]), .B1(N96), 
        .Y(N987) );
  AOI22X1TF U590 ( .A0(SUM_AB[6]), .A1(N171), .B0(N991), .B1(N1014), .Y(N992)
         );
  AOI22X1TF U591 ( .A0(DIVISION_HEAD[6]), .A1(N69), .B0(ZTEMP[6]), .B1(N96), 
        .Y(N993) );
  AOI22X1TF U592 ( .A0(SUM_AB[2]), .A1(N171), .B0(N979), .B1(N1014), .Y(N980)
         );
  AOI22X1TF U593 ( .A0(DIVISION_HEAD[2]), .A1(N69), .B0(ZTEMP[2]), .B1(N96), 
        .Y(N981) );
  AOI22X1TF U594 ( .A0(SUM_AB[1]), .A1(N171), .B0(N976), .B1(N1014), .Y(N977)
         );
  AOI22X1TF U595 ( .A0(DIVISION_HEAD[1]), .A1(N69), .B0(ZTEMP[1]), .B1(N96), 
        .Y(N978) );
  OAI211X1TF U596 ( .A0(N75), .A1(N369), .B0(N644), .C0(N368), .Y(N721) );
  AOI22X1TF U597 ( .A0(STEP[3]), .A1(N641), .B0(N375), .B1(N573), .Y(N368) );
  OAI211X1TF U598 ( .A0(N155), .A1(N941), .B0(N843), .C0(N842), .Y(N679) );
  AOI211X1TF U599 ( .A0(OPER_A[3]), .A1(N841), .B0(N840), .C0(N839), .Y(N842)
         );
  OAI31X1TF U600 ( .A0(N931), .A1(N838), .A2(OPER_A[3]), .B0(N187), .Y(N839)
         );
  AOI21X1TF U601 ( .A0(C152_DATA4_3), .A1(N200), .B0(N895), .Y(N187) );
  OAI32X1TF U602 ( .A0(N163), .A1(N934), .A2(N837), .B0(N932), .B1(N163), .Y(
        N840) );
  OAI21X1TF U603 ( .A0(N931), .A1(N836), .B0(N929), .Y(N841) );
  AOI31X1TF U604 ( .A0(N898), .A1(N163), .A2(N837), .B0(N871), .Y(N843) );
  OAI22X1TF U605 ( .A0(N514), .A1(N513), .B0(N512), .B1(N133), .Y(N708) );
  OAI21X1TF U606 ( .A0(N507), .A1(N1008), .B0(N506), .Y(N508) );
  AOI211X1TF U607 ( .A0(SUM_AB[11]), .A1(N84), .B0(N505), .C0(N504), .Y(N506)
         );
  OAI22X1TF U608 ( .A0(N136), .A1(N734), .B0(N501), .B1(N59), .Y(N505) );
  AOI22X1TF U609 ( .A0(N476), .A1(N131), .B0(N442), .B1(N461), .Y(N714) );
  AOI21X1TF U610 ( .A0(DIVISION_HEAD[8]), .A1(N79), .B0(N435), .Y(N436) );
  OAI22X1TF U611 ( .A0(N131), .A1(N455), .B0(N507), .B1(N990), .Y(N435) );
  AOI22X1TF U612 ( .A0(DIVISION_HEAD[10]), .A1(N99), .B0(X_IN[10]), .B1(N62), 
        .Y(N438) );
  OAI22X1TF U613 ( .A0(N443), .A1(N608), .B0(N558), .B1(N477), .Y(N441) );
  AOI32X1TF U614 ( .A0(N403), .A1(N461), .A2(N402), .B0(N476), .B1(N119), .Y(
        N718) );
  AOI211X1TF U615 ( .A0(N494), .A1(N976), .B0(N401), .C0(N400), .Y(N402) );
  OAI211X1TF U616 ( .A0(N558), .A1(N433), .B0(N399), .C0(N398), .Y(N400) );
  AOI21X1TF U617 ( .A0(DIVISION_HEAD[4]), .A1(N80), .B0(N397), .Y(N398) );
  OAI22X1TF U618 ( .A0(N119), .A1(N455), .B0(N747), .B1(N608), .Y(N397) );
  OAI22X1TF U619 ( .A0(N464), .A1(N396), .B0(N489), .B1(N805), .Y(N401) );
  AOI21X1TF U620 ( .A0(SUM_AB[1]), .A1(SUM_AB[0]), .B0(N405), .Y(N976) );
  AOI32X1TF U621 ( .A0(N462), .A1(N461), .A2(N460), .B0(N476), .B1(N127), .Y(
        N712) );
  OAI211X1TF U622 ( .A0(N507), .A1(N996), .B0(N457), .C0(N456), .Y(N458) );
  AOI22X1TF U623 ( .A0(DIVISION_HEAD[12]), .A1(N99), .B0(X_IN[12]), .B1(N62), 
        .Y(N456) );
  AOI22X1TF U624 ( .A0(DIVISION_HEAD[11]), .A1(N804), .B0(DIVISION_HEAD[10]), 
        .B1(N79), .Y(N457) );
  OAI22X1TF U625 ( .A0(N464), .A1(N608), .B0(N558), .B1(N499), .Y(N459) );
  AOI32X1TF U626 ( .A0(N423), .A1(N461), .A2(N422), .B0(N476), .B1(N42), .Y(
        N716) );
  AOI211X1TF U627 ( .A0(DIVISION_HEAD[8]), .A1(N99), .B0(N421), .C0(N420), .Y(
        N422) );
  OAI211X1TF U628 ( .A0(N558), .A1(N453), .B0(N419), .C0(N418), .Y(N420) );
  AOI21X1TF U629 ( .A0(DIVISION_HEAD[6]), .A1(N80), .B0(N417), .Y(N418) );
  OAI22X1TF U630 ( .A0(N42), .A1(N455), .B0(N507), .B1(N984), .Y(N417) );
  INVX2TF U631 ( .A(N494), .Y(N507) );
  AOI22X1TF U632 ( .A0(N174), .A1(N445), .B0(X_IN[1]), .B1(N800), .Y(N419) );
  OAI21X1TF U633 ( .A0(N503), .A1(N805), .B0(N414), .Y(N421) );
  AOI22X1TF U634 ( .A0(X_IN[8]), .A1(N63), .B0(X_IN[9]), .B1(N67), .Y(N414) );
  OAI211X1TF U635 ( .A0(N852), .A1(N851), .B0(N850), .C0(N849), .Y(N678) );
  AOI32X1TF U636 ( .A0(N898), .A1(OPER_B[4]), .A2(N848), .B0(N873), .B1(
        OPER_B[4]), .Y(N849) );
  AOI211X1TF U637 ( .A0(N853), .A1(OPER_B[5]), .B0(N847), .C0(N846), .Y(N850)
         );
  OAI31X1TF U638 ( .A0(N931), .A1(N845), .A2(OPER_A[4]), .B0(N188), .Y(N846)
         );
  AOI21X1TF U639 ( .A0(N200), .A1(C152_DATA4_4), .B0(N189), .Y(N188) );
  NOR3X1TF U640 ( .A(OPER_B[4]), .B(N848), .C(N934), .Y(N847) );
  AOI21X1TF U641 ( .A0(N928), .A1(N845), .B0(N844), .Y(N851) );
  OAI211X1TF U642 ( .A0(N161), .A1(N614), .B0(N630), .C0(N613), .Y(N700) );
  AOI21X1TF U643 ( .A0(N641), .A1(N147), .B0(N612), .Y(N613) );
  NOR3X1TF U644 ( .A(STEP[3]), .B(N75), .C(N603), .Y(N947) );
  AOI211X1TF U645 ( .A0(N822), .A1(N375), .B0(N372), .C0(N371), .Y(N611) );
  AOI21X1TF U646 ( .A0(N385), .A1(N370), .B0(N774), .Y(N371) );
  NOR2X1TF U647 ( .A(N73), .B(N821), .Y(N375) );
  OAI211X1TF U648 ( .A0(N645), .A1(N134), .B0(N644), .C0(N643), .Y(N696) );
  NOR2X1TF U649 ( .A(N648), .B(N362), .Y(N644) );
  INVX2TF U650 ( .A(N649), .Y(N648) );
  AOI21X1TF U651 ( .A0(N642), .A1(N944), .B0(N641), .Y(N645) );
  NOR4BX1TF U652 ( .AN(N345), .B(N926), .C(N347), .D(N819), .Y(N201) );
  OAI31X1TF U653 ( .A0(OPER_B[12]), .A1(N339), .A2(N934), .B0(N823), .Y(N347)
         );
  NOR2X1TF U654 ( .A(OPER_B[11]), .B(N933), .Y(N339) );
  AOI32X1TF U655 ( .A0(N944), .A1(OPER_B[12]), .A2(N344), .B0(N203), .B1(
        OPER_B[12]), .Y(N345) );
  OAI31X1TF U656 ( .A0(N907), .A1(OPER_B[11]), .A2(N933), .B0(N857), .Y(N344)
         );
  INVX2TF U657 ( .A(N918), .Y(N907) );
  AOI22X1TF U658 ( .A0(N341), .A1(N928), .B0(OPER_A[12]), .B1(N844), .Y(N346)
         );
  NOR2X1TF U659 ( .A(N930), .B(OPER_A[11]), .Y(N340) );
  INVX2TF U660 ( .A(OPER_A[8]), .Y(N885) );
  INVX2TF U661 ( .A(OPER_A[10]), .Y(N911) );
  OAI21X1TF U662 ( .A0(N82), .A1(N548), .B0(N94), .Y(C2_Z_12) );
  OAI22X1TF U663 ( .A0(N81), .A1(N759), .B0(N185), .B1(OFFSET[6]), .Y(C2_Z_8)
         );
  OAI22X1TF U664 ( .A0(N82), .A1(N781), .B0(N94), .B1(OFFSET[7]), .Y(C2_Z_9)
         );
  OAI22X1TF U665 ( .A0(N81), .A1(N547), .B0(N185), .B1(OFFSET[8]), .Y(C2_Z_10)
         );
  OAI22X1TF U666 ( .A0(N81), .A1(N803), .B0(N185), .B1(OFFSET[9]), .Y(C2_Z_11)
         );
  AOI32X1TF U667 ( .A0(N820), .A1(N944), .A2(N821), .B0(N637), .B1(N944), .Y(
        N643) );
  OAI22X1TF U668 ( .A0(N120), .A1(N952), .B0(N821), .B1(N965), .Y(N637) );
  AOI211X1TF U669 ( .A0(N641), .A1(N120), .B0(N636), .C0(N635), .Y(N640) );
  AOI21X1TF U670 ( .A0(DP_OP_333_124_4748_N43), .A1(N602), .B0(N601), .Y(N630)
         );
  OAI21X1TF U671 ( .A0(N600), .A1(N599), .B0(N598), .Y(N601) );
  OR2X2TF U672 ( .A(N828), .B(N830), .Y(N194) );
  AOI21X1TF U673 ( .A0(N928), .A1(N829), .B0(N844), .Y(N828) );
  AOI21X1TF U674 ( .A0(N88), .A1(C152_DATA4_1), .B0(N874), .Y(N195) );
  AOI211X1TF U675 ( .A0(N853), .A1(OPER_B[2]), .B0(N826), .C0(N825), .Y(N827)
         );
  NOR3X1TF U676 ( .A(N829), .B(OPER_A[1]), .C(N931), .Y(N825) );
  OAI32X1TF U677 ( .A0(N162), .A1(OPER_B[0]), .A2(N934), .B0(N932), .B1(N162), 
        .Y(N826) );
  INVX2TF U678 ( .A(N882), .Y(N853) );
  OAI31X1TF U679 ( .A0(OPER_B[1]), .A1(N89), .A2(N164), .B0(N823), .Y(N824) );
  OAI21X1TF U680 ( .A0(N451), .A1(N450), .B0(N461), .Y(N452) );
  AOI22X1TF U681 ( .A0(DIVISION_HEAD[11]), .A1(N99), .B0(X_IN[12]), .B1(N67), 
        .Y(N446) );
  AOI22X1TF U682 ( .A0(N61), .A1(N445), .B0(X_IN[11]), .B1(N63), .Y(N447) );
  AOI22X1TF U683 ( .A0(SUM_AB[6]), .A1(N85), .B0(N494), .B1(N991), .Y(N448) );
  AOI21X1TF U684 ( .A0(SUM_AB[6]), .A1(N444), .B0(N454), .Y(N991) );
  AOI22X1TF U685 ( .A0(XTEMP[11]), .A1(N80), .B0(X_IN[11]), .B1(N445), .Y(N354) );
  OAI211X1TF U686 ( .A0(N882), .A1(N139), .B0(N881), .C0(N880), .Y(N675) );
  AOI211X1TF U687 ( .A0(OPER_A[7]), .A1(N878), .B0(N877), .C0(N876), .Y(N881)
         );
  AOI211X1TF U688 ( .A0(N45), .A1(N963), .B0(SIGN_Y), .C0(N906), .Y(N926) );
  OAI21X1TF U689 ( .A0(N82), .A1(N184), .B0(N94), .Y(C2_Z_1) );
  INVX2TF U690 ( .A(Y_IN[1]), .Y(N184) );
  OAI22X1TF U691 ( .A0(N82), .A1(N183), .B0(N94), .B1(OFFSET[1]), .Y(C2_Z_3)
         );
  INVX2TF U692 ( .A(Y_IN[3]), .Y(N183) );
  OAI22X1TF U693 ( .A0(N81), .A1(N182), .B0(N185), .B1(OFFSET[2]), .Y(C2_Z_4)
         );
  INVX2TF U694 ( .A(Y_IN[4]), .Y(N182) );
  OAI22X1TF U695 ( .A0(N82), .A1(N181), .B0(N94), .B1(OFFSET[3]), .Y(C2_Z_5)
         );
  INVX2TF U696 ( .A(N172), .Y(N181) );
  OAI22X1TF U697 ( .A0(N82), .A1(N173), .B0(N94), .B1(OFFSET[5]), .Y(C2_Z_7)
         );
  INVX2TF U698 ( .A(N932), .Y(N873) );
  INVX2TF U699 ( .A(N862), .Y(N858) );
  INVX2TF U700 ( .A(N934), .Y(N898) );
  OAI21X1TF U701 ( .A0(N931), .A1(N879), .B0(N929), .Y(N878) );
  INVX2TF U702 ( .A(N838), .Y(N836) );
  INVX2TF U703 ( .A(OPER_A[4]), .Y(N852) );
  INVX2TF U704 ( .A(OPER_A[6]), .Y(N864) );
  AOI32X1TF U705 ( .A0(N432), .A1(N461), .A2(N431), .B0(N476), .B1(N130), .Y(
        N715) );
  AOI211X1TF U706 ( .A0(N494), .A1(N985), .B0(N430), .C0(N429), .Y(N431) );
  AOI22X1TF U707 ( .A0(N174), .A1(N800), .B0(N56), .B1(N445), .Y(N426) );
  AOI22X1TF U708 ( .A0(DIVISION_HEAD[9]), .A1(N99), .B0(X_IN[9]), .B1(N62), 
        .Y(N427) );
  AOI22X1TF U709 ( .A0(X_IN[10]), .A1(N66), .B0(X_IN[11]), .B1(N83), .Y(N428)
         );
  AOI21X1TF U710 ( .A0(SUM_AB[4]), .A1(N424), .B0(N434), .Y(N985) );
  OAI21X1TF U711 ( .A0(N758), .A1(N146), .B0(N757), .Y(N687) );
  OAI21X1TF U712 ( .A0(N756), .A1(N755), .B0(N777), .Y(N757) );
  OAI211X1TF U713 ( .A0(N144), .A1(N774), .B0(N754), .C0(N753), .Y(N755) );
  AOI22X1TF U714 ( .A0(DIVISION_REMA[6]), .A1(N80), .B0(SUM_AB[7]), .B1(N797), 
        .Y(N753) );
  OAI211X1TF U715 ( .A0(N808), .A1(N996), .B0(N752), .C0(N751), .Y(N756) );
  AOI22X1TF U716 ( .A0(X_IN[1]), .A1(N83), .B0(X_IN[0]), .B1(N67), .Y(N751) );
  AOI32X1TF U717 ( .A0(N1018), .A1(N975), .A2(N1009), .B0(N974), .B1(N975), 
        .Y(N669) );
  INVX2TF U718 ( .A(SUM_AB[0]), .Y(N974) );
  AOI22X1TF U719 ( .A0(DIVISION_HEAD[0]), .A1(N68), .B0(ZTEMP[0]), .B1(N1010), 
        .Y(N975) );
  AOI22X1TF U720 ( .A0(N170), .A1(N144), .B0(N778), .B1(N777), .Y(N686) );
  INVX2TF U721 ( .A(N170), .Y(N777) );
  AOI211X1TF U722 ( .A0(DIVISION_REMA[7]), .A1(N80), .B0(N776), .C0(N775), .Y(
        N778) );
  OAI211X1TF U723 ( .A0(N148), .A1(N774), .B0(N773), .C0(N772), .Y(N775) );
  AOI22X1TF U724 ( .A0(N771), .A1(N770), .B0(N997), .B1(N794), .Y(N772) );
  AOI32X1TF U725 ( .A0(N769), .A1(N768), .A2(N767), .B0(N766), .B1(N768), .Y(
        N770) );
  INVX2TF U726 ( .A(N174), .Y(N769) );
  AOI22X1TF U727 ( .A0(DIVISION_REMA[8]), .A1(N760), .B0(SUM_AB[8]), .B1(N797), 
        .Y(N773) );
  OAI31X1TF U728 ( .A0(N629), .A1(N628), .A2(N627), .B0(N626), .Y(N698) );
  AOI22X1TF U729 ( .A0(\INDEX[2] ), .A1(N625), .B0(N624), .B1(N623), .Y(N626)
         );
  OAI21X1TF U730 ( .A0(N622), .A1(N628), .B0(N621), .Y(N625) );
  OAI211X1TF U731 ( .A0(N1009), .A1(N1008), .B0(N1007), .C0(N1006), .Y(N658)
         );
  AOI22X1TF U732 ( .A0(DIVISION_HEAD[11]), .A1(N69), .B0(ZTEMP[11]), .B1(N1010), .Y(N1007) );
  OAI211X1TF U733 ( .A0(N1009), .A1(N996), .B0(N995), .C0(N994), .Y(N662) );
  AOI22X1TF U734 ( .A0(DIVISION_HEAD[7]), .A1(N68), .B0(ZTEMP[7]), .B1(N1010), 
        .Y(N995) );
  OAI21X1TF U735 ( .A0(N454), .A1(N453), .B0(N463), .Y(N996) );
  OAI211X1TF U736 ( .A0(N1009), .A1(N1002), .B0(N1001), .C0(N1000), .Y(N660)
         );
  AOI22X1TF U737 ( .A0(DIVISION_HEAD[9]), .A1(N68), .B0(ZTEMP[9]), .B1(N1010), 
        .Y(N1001) );
  OAI211X1TF U738 ( .A0(N1009), .A1(N990), .B0(N989), .C0(N988), .Y(N664) );
  AOI22X1TF U739 ( .A0(DIVISION_HEAD[5]), .A1(N68), .B0(ZTEMP[5]), .B1(N1010), 
        .Y(N989) );
  OAI211X1TF U740 ( .A0(N1009), .A1(N984), .B0(N983), .C0(N982), .Y(N666) );
  NOR3X1TF U741 ( .A(N64), .B(N157), .C(N963), .Y(N962) );
  AOI22X1TF U742 ( .A0(DIVISION_HEAD[3]), .A1(N68), .B0(ZTEMP[3]), .B1(N1010), 
        .Y(N983) );
  AOI211X4TF U743 ( .A0(N973), .A1(N972), .B0(N971), .C0(N1010), .Y(N1014) );
  AOI31X1TF U744 ( .A0(N958), .A1(N957), .A2(N956), .B0(N955), .Y(N961) );
  OAI31X1TF U745 ( .A0(N954), .A1(N953), .A2(N952), .B0(N951), .Y(N955) );
  INVX2TF U746 ( .A(N968), .Y(N971) );
  NOR2X1TF U747 ( .A(N629), .B(N623), .Y(N621) );
  AOI21X1TF U748 ( .A0(\INDEX[2] ), .A1(N624), .B0(N376), .Y(N623) );
  INVX2TF U749 ( .A(N619), .Y(N629) );
  INVX2TF U750 ( .A(N247), .Y(N633) );
  AOI31X1TF U751 ( .A0(N954), .A1(N370), .A2(N385), .B0(N774), .Y(N247) );
  OAI21X1TF U752 ( .A0(N351), .A1(N246), .B0(N78), .Y(N361) );
  INVX2TF U753 ( .A(N616), .Y(N624) );
  NOR2X1TF U754 ( .A(N965), .B(N832), .Y(N859) );
  AOI221X1TF U755 ( .A0(N128), .A1(N138), .B0(N160), .B1(N91), .C0(N817), .Y(
        N818) );
  AOI22X1TF U756 ( .A0(\INDEX[2] ), .A1(N90), .B0(N124), .B1(\RSHT_BITS[3] ), 
        .Y(N816) );
  NOR3X1TF U757 ( .A(N64), .B(N906), .C(N970), .Y(N819) );
  AOI21X2TF U758 ( .A0(N78), .A1(N917), .B0(N203), .Y(N932) );
  INVX2TF U759 ( .A(N857), .Y(N917) );
  AOI32X1TF U760 ( .A0(N605), .A1(N343), .A2(N822), .B0(N948), .B1(N342), .Y(
        N857) );
  INVX2TF U761 ( .A(N943), .Y(N948) );
  AND2X2TF U762 ( .A(N925), .B(N186), .Y(N200) );
  NAND2X2TF U763 ( .A(N564), .B(N343), .Y(N912) );
  INVX2TF U764 ( .A(N342), .Y(N343) );
  INVX2TF U765 ( .A(N929), .Y(N844) );
  NAND2X2TF U766 ( .A(N908), .B(N892), .Y(N929) );
  INVX2TF U767 ( .A(N833), .Y(N908) );
  AOI21X1TF U768 ( .A0(N564), .A1(N342), .B0(N563), .Y(N833) );
  INVX2TF U769 ( .A(N338), .Y(N957) );
  INVX2TF U770 ( .A(N565), .Y(N950) );
  AOI21X1TF U771 ( .A0(N822), .A1(N821), .B0(N820), .Y(N831) );
  NOR2X2TF U772 ( .A(N603), .B(N631), .Y(N822) );
  AOI32X1TF U773 ( .A0(N943), .A1(N951), .A2(N369), .B0(N953), .B1(N951), .Y(
        N336) );
  INVX2TF U774 ( .A(N603), .Y(N642) );
  OAI21X1TF U775 ( .A0(N338), .A1(N942), .B0(N334), .Y(N607) );
  OAI21X1TF U776 ( .A0(N570), .A1(N564), .B0(N335), .Y(N334) );
  INVX2TF U777 ( .A(N820), .Y(N378) );
  OAI31X1TF U778 ( .A0(N328), .A1(DIVISION_HEAD[10]), .A2(N547), .B0(N327), 
        .Y(N329) );
  AOI22X1TF U779 ( .A0(Y_IN[11]), .A1(N127), .B0(N326), .B1(N325), .Y(N327) );
  OAI22X1TF U780 ( .A0(DIVISION_HEAD[8]), .A1(N759), .B0(DIVISION_HEAD[9]), 
        .B1(N781), .Y(N325) );
  INVX2TF U781 ( .A(N324), .Y(N326) );
  NOR2X1TF U782 ( .A(Y_IN[11]), .B(N127), .Y(N328) );
  AOI22X1TF U783 ( .A0(DIVISION_HEAD[10]), .A1(N547), .B0(DIVISION_HEAD[9]), 
        .B1(N781), .Y(N322) );
  NOR2X1TF U784 ( .A(N57), .B(N42), .Y(N319) );
  AOI32X1TF U785 ( .A0(N796), .A1(N814), .A2(N795), .B0(N812), .B1(N150), .Y(
        N684) );
  AOI21X1TF U786 ( .A0(N794), .A1(N1003), .B0(N793), .Y(N795) );
  AOI22X1TF U787 ( .A0(N174), .A1(N63), .B0(N175), .B1(N83), .Y(N789) );
  AOI22X1TF U788 ( .A0(DIVISION_HEAD[0]), .A1(N79), .B0(DIVISION_HEAD[1]), 
        .B1(N804), .Y(N790) );
  AOI22X1TF U789 ( .A0(Y_IN[10]), .A1(N788), .B0(N56), .B1(N67), .Y(N791) );
  AOI21X1TF U790 ( .A0(SUM_AB[10]), .A1(N487), .B0(N500), .Y(N1003) );
  AOI22X1TF U791 ( .A0(N798), .A1(SUM_AB[1]), .B0(SUM_AB[10]), .B1(N98), .Y(
        N796) );
  OAI21X1TF U792 ( .A0(N812), .A1(N555), .B0(N554), .Y(N706) );
  OAI21X1TF U793 ( .A0(N812), .A1(N804), .B0(DIVISION_HEAD[3]), .Y(N554) );
  AOI211X1TF U794 ( .A0(DIVISION_HEAD[2]), .A1(N80), .B0(N553), .C0(N552), .Y(
        N555) );
  AOI22X1TF U795 ( .A0(N798), .A1(SUM_AB[3]), .B0(N1012), .B1(N794), .Y(N549)
         );
  AOI22X1TF U796 ( .A0(N944), .A1(SUM_AB[12]), .B0(N61), .B1(N67), .Y(N550) );
  AOI22X1TF U797 ( .A0(N175), .A1(N63), .B0(X_IN[6]), .B1(N83), .Y(N551) );
  OAI22X1TF U798 ( .A0(N548), .A1(N802), .B0(N547), .B1(N59), .Y(N553) );
  INVX2TF U799 ( .A(Y_IN[12]), .Y(N548) );
  AOI32X1TF U800 ( .A0(N394), .A1(N393), .A2(N392), .B0(N476), .B1(N393), .Y(
        N719) );
  OAI211X1TF U801 ( .A0(N390), .A1(N558), .B0(N389), .C0(N388), .Y(N391) );
  AOI22X1TF U802 ( .A0(X_IN[6]), .A1(N67), .B0(N61), .B1(N63), .Y(N388) );
  AOI22X1TF U803 ( .A0(DIVISION_HEAD[5]), .A1(N99), .B0(N176), .B1(N83), .Y(
        N389) );
  AOI22X1TF U804 ( .A0(DIVISION_HEAD[3]), .A1(N80), .B0(SUM_AB[0]), .B1(N382), 
        .Y(N394) );
  OAI22X1TF U805 ( .A0(N476), .A1(N475), .B0(N474), .B1(N135), .Y(N711) );
  NAND2X2TF U806 ( .A(N455), .B(N461), .Y(N472) );
  AOI211X1TF U807 ( .A0(N997), .A1(N494), .B0(N471), .C0(N470), .Y(N475) );
  OAI211X1TF U808 ( .A0(N469), .A1(N608), .B0(N468), .C0(N467), .Y(N470) );
  AOI22X1TF U809 ( .A0(XTEMP[9]), .A1(N99), .B0(N798), .B1(SUM_AB[12]), .Y(
        N467) );
  NOR2X1TF U810 ( .A(DIVISION_HEAD[12]), .B(N473), .Y(N466) );
  AOI22X1TF U811 ( .A0(X_IN[8]), .A1(N465), .B0(INTADD_0_N1), .B1(N489), .Y(
        N473) );
  INVX2TF U812 ( .A(INTADD_0_N1), .Y(N465) );
  OAI22X1TF U813 ( .A0(N127), .A1(N47), .B0(N464), .B1(N59), .Y(N471) );
  OAI22X1TF U814 ( .A0(N170), .A1(N743), .B0(N758), .B1(N145), .Y(N689) );
  AOI211X1TF U815 ( .A0(SUM_AB[5]), .A1(N98), .B0(N742), .C0(N741), .Y(N743)
         );
  OAI211X1TF U816 ( .A0(N808), .A1(N990), .B0(N754), .C0(N740), .Y(N741) );
  OAI21X1TF U817 ( .A0(N434), .A1(N433), .B0(N444), .Y(N990) );
  INVX2TF U818 ( .A(N802), .Y(N788) );
  OAI22X1TF U819 ( .A0(N170), .A1(N733), .B0(N758), .B1(N143), .Y(N691) );
  AOI211X1TF U820 ( .A0(SUM_AB[3]), .A1(N98), .B0(N732), .C0(N731), .Y(N733)
         );
  OAI211X1TF U821 ( .A0(N808), .A1(N984), .B0(N754), .C0(N730), .Y(N731) );
  AOI222X4TF U822 ( .A0(N764), .A1(N62), .B0(N762), .B1(N66), .C0(N557), .C1(
        N83), .Y(N754) );
  OAI21X1TF U823 ( .A0(N416), .A1(N415), .B0(N424), .Y(N984) );
  OAI22X1TF U824 ( .A0(N729), .A1(N802), .B0(N153), .B1(N734), .Y(N732) );
  AOI32X1TF U825 ( .A0(N413), .A1(N461), .A2(N412), .B0(N476), .B1(N126), .Y(
        N717) );
  AOI211X1TF U826 ( .A0(DIVISION_HEAD[7]), .A1(N99), .B0(N411), .C0(N410), .Y(
        N412) );
  OAI211X1TF U827 ( .A0(N59), .A1(N747), .B0(N409), .C0(N408), .Y(N410) );
  AOI21X1TF U828 ( .A0(N494), .A1(N979), .B0(N407), .Y(N408) );
  AOI21X1TF U829 ( .A0(SUM_AB[2]), .A1(N406), .B0(N416), .Y(N979) );
  NOR2X1TF U830 ( .A(SUM_AB[0]), .B(SUM_AB[1]), .Y(N405) );
  NOR2X2TF U831 ( .A(N395), .B(N1017), .Y(N494) );
  AOI22X1TF U832 ( .A0(X_IN[1]), .A1(N445), .B0(N798), .B1(SUM_AB[6]), .Y(N409) );
  INVX2TF U833 ( .A(N608), .Y(N445) );
  NAND2X2TF U834 ( .A(MODE_TYPE[1]), .B(N353), .Y(N608) );
  OAI21X1TF U835 ( .A0(N501), .A1(N805), .B0(N404), .Y(N411) );
  AOI22X1TF U836 ( .A0(X_IN[8]), .A1(N67), .B0(N176), .B1(N63), .Y(N404) );
  OAI211X1TF U837 ( .A0(N64), .A1(N376), .B0(N360), .C0(N349), .Y(N350) );
  NOR2X1TF U838 ( .A(N372), .B(N946), .Y(N360) );
  INVX2TF U839 ( .A(N395), .Y(N372) );
  INVX2TF U840 ( .A(N617), .Y(N376) );
  NOR2X1TF U841 ( .A(N125), .B(N747), .Y(INTADD_0_CI) );
  INVX2TF U842 ( .A(N605), .Y(N821) );
  NOR2X1TF U843 ( .A(PRE_WORK), .B(N365), .Y(N602) );
  AOI32X1TF U844 ( .A0(N787), .A1(N814), .A2(N786), .B0(N812), .B1(N148), .Y(
        N685) );
  OAI211X1TF U845 ( .A0(N808), .A1(N1002), .B0(N783), .C0(N782), .Y(N784) );
  AOI22X1TF U846 ( .A0(DIVISION_HEAD[1]), .A1(N77), .B0(X_IN[1]), .B1(N62), 
        .Y(N782) );
  OAI21X1TF U847 ( .A0(N478), .A1(N477), .B0(N487), .Y(N1002) );
  OAI21X1TF U848 ( .A0(N781), .A1(N802), .B0(N780), .Y(N785) );
  AOI22X1TF U849 ( .A0(DIVISION_REMA[8]), .A1(N79), .B0(N798), .B1(SUM_AB[0]), 
        .Y(N780) );
  AOI22X1TF U850 ( .A0(DIVISION_HEAD[0]), .A1(N804), .B0(SUM_AB[9]), .B1(N98), 
        .Y(N787) );
  NOR2X1TF U851 ( .A(N332), .B(N370), .Y(ALU_IS_DONE) );
  OAI211X1TF U852 ( .A0(N126), .A1(N54), .B0(N208), .C0(N207), .Y(FOUT[0]) );
  AOI32X1TF U853 ( .A0(N815), .A1(N814), .A2(N813), .B0(N812), .B1(N43), .Y(
        N683) );
  AOI211X1TF U854 ( .A0(DIVISION_HEAD[3]), .A1(N76), .B0(N810), .C0(N809), .Y(
        N813) );
  OAI211X1TF U855 ( .A0(N808), .A1(N1008), .B0(N807), .C0(N806), .Y(N809) );
  AOI22X1TF U856 ( .A0(N56), .A1(N62), .B0(N61), .B1(N83), .Y(N806) );
  AND2X2TF U857 ( .A(N761), .B(N766), .Y(N763) );
  INVX2TF U858 ( .A(N387), .Y(N771) );
  AOI22X1TF U859 ( .A0(DIVISION_HEAD[1]), .A1(N79), .B0(DIVISION_HEAD[2]), 
        .B1(N804), .Y(N807) );
  INVX2TF U860 ( .A(N455), .Y(N804) );
  OAI21X1TF U861 ( .A0(N500), .A1(N499), .B0(N1013), .Y(N1008) );
  INVX2TF U862 ( .A(SUM_AB[11]), .Y(N499) );
  INVX2TF U863 ( .A(SUM_AB[9]), .Y(N477) );
  INVX2TF U864 ( .A(SUM_AB[7]), .Y(N453) );
  INVX2TF U865 ( .A(SUM_AB[5]), .Y(N433) );
  INVX2TF U866 ( .A(SUM_AB[3]), .Y(N415) );
  INVX2TF U867 ( .A(N794), .Y(N808) );
  NOR2X2TF U868 ( .A(N1017), .B(N649), .Y(N794) );
  INVX2TF U869 ( .A(SUM_AB[12]), .Y(N1017) );
  OAI21X1TF U870 ( .A0(N803), .A1(N802), .B0(N801), .Y(N810) );
  INVX2TF U871 ( .A(N812), .Y(N814) );
  NOR3X2TF U872 ( .A(N73), .B(N604), .C(N631), .Y(N617) );
  AND2X2TF U873 ( .A(N646), .B(N639), .Y(N545) );
  INVX2TF U874 ( .A(N353), .Y(N639) );
  INVX2TF U875 ( .A(N301), .Y(N762) );
  OAI211X1TF U876 ( .A0(X_IN[12]), .A1(N547), .B0(N300), .C0(N299), .Y(N301)
         );
  OAI22X1TF U877 ( .A0(Y_IN[10]), .A1(N298), .B0(N297), .B1(N296), .Y(N299) );
  OAI22X1TF U878 ( .A0(X_IN[10]), .A1(N295), .B0(N86), .B1(N781), .Y(N296) );
  OAI21X1TF U879 ( .A0(Y_IN[9]), .A1(N177), .B0(Y_IN[8]), .Y(N295) );
  NOR2X1TF U880 ( .A(N57), .B(N501), .Y(N290) );
  OAI22X1TF U881 ( .A0(N175), .A1(N736), .B0(X_IN[5]), .B1(N729), .Y(N285) );
  INVX2TF U882 ( .A(N176), .Y(N469) );
  INVX2TF U883 ( .A(X_IN[9]), .Y(N501) );
  NOR2X1TF U884 ( .A(Y_IN[9]), .B(N177), .Y(N294) );
  NOR2X1TF U885 ( .A(Y_IN[12]), .B(Y_IN[11]), .Y(N300) );
  NOR2X1TF U886 ( .A(Y_IN[9]), .B(N298), .Y(N280) );
  NOR2X1TF U887 ( .A(N57), .B(N503), .Y(N276) );
  OAI22X1TF U888 ( .A0(X_IN[6]), .A1(N729), .B0(X_IN[5]), .B1(N736), .Y(N271)
         );
  OR2X2TF U889 ( .A(MODE_TYPE[0]), .B(N306), .Y(N766) );
  INVX2TF U890 ( .A(MODE_TYPE[1]), .Y(N306) );
  OAI31X1TF U891 ( .A0(N268), .A1(N86), .A2(N547), .B0(N267), .Y(N269) );
  OAI31X1TF U892 ( .A0(N266), .A1(N265), .A2(N264), .B0(N263), .Y(N267) );
  AOI22X1TF U893 ( .A0(N86), .A1(N547), .B0(X_IN[12]), .B1(N803), .Y(N263) );
  INVX2TF U894 ( .A(Y_IN[11]), .Y(N803) );
  NOR2X1TF U895 ( .A(X_IN[10]), .B(N781), .Y(N264) );
  AOI211X1TF U896 ( .A0(X_IN[10]), .A1(N781), .B0(X_IN[9]), .C0(N759), .Y(N265) );
  NOR2X1TF U897 ( .A(N57), .B(N489), .Y(N258) );
  NOR2X1TF U898 ( .A(N172), .B(N464), .Y(N254) );
  AOI211X1TF U899 ( .A0(N175), .A1(N729), .B0(N56), .C0(N736), .Y(N251) );
  AOI22X1TF U900 ( .A0(X_IN[3]), .A1(N736), .B0(N174), .B1(N308), .Y(N249) );
  INVX2TF U901 ( .A(X_IN[6]), .Y(N464) );
  NOR2X1TF U902 ( .A(Y_IN[9]), .B(N503), .Y(N262) );
  NOR2X1TF U903 ( .A(Y_IN[11]), .B(N298), .Y(N268) );
  INVX2TF U904 ( .A(X_IN[12]), .Y(N298) );
  INVX2TF U905 ( .A(N332), .Y(N385) );
  AOI22X1TF U906 ( .A0(N798), .A1(SUM_AB[2]), .B0(SUM_AB[11]), .B1(N98), .Y(
        N815) );
  INVX2TF U907 ( .A(N305), .Y(N627) );
  OAI21X1TF U908 ( .A0(N44), .A1(N70), .B0(N242), .Y(OPER_A[12]) );
  OAI21X1TF U909 ( .A0(N130), .A1(N70), .B0(N233), .Y(OPER_A[4]) );
  OAI21X1TF U910 ( .A0(N132), .A1(N70), .B0(N235), .Y(OPER_A[6]) );
  OAI21X1TF U911 ( .A0(N127), .A1(N48), .B0(N236), .Y(OPER_A[7]) );
  OAI21X1TF U912 ( .A0(N135), .A1(N70), .B0(N237), .Y(OPER_A[8]) );
  OAI21X1TF U913 ( .A0(N48), .A1(N39), .B0(N238), .Y(OPER_A[9]) );
  OAI21X1TF U914 ( .A0(N70), .A1(N136), .B0(N239), .Y(OPER_A[10]) );
  OAI21X1TF U915 ( .A0(N48), .A1(N133), .B0(N240), .Y(OPER_A[11]) );
  INVX2TF U916 ( .A(N558), .Y(N798) );
  AOI31X1TF U917 ( .A0(N509), .A1(N136), .A2(N495), .B0(N490), .Y(N491) );
  AOI31X1TF U918 ( .A0(N95), .A1(N133), .A2(N510), .B0(N508), .Y(N513) );
  AOI22X1TF U919 ( .A0(N509), .A1(\INTADD_0_SUM[5] ), .B0(N798), .B1(
        SUM_AB[10]), .Y(N449) );
  AOI21X1TF U920 ( .A0(N95), .A1(N357), .B0(N514), .Y(N358) );
  INVX2TF U921 ( .A(N1010), .Y(N967) );
  AOI31X1TF U922 ( .A0(X_IN[0]), .A1(N95), .A2(N125), .B0(N391), .Y(N392) );
  AOI21X1TF U923 ( .A0(N95), .A1(N473), .B0(N472), .Y(N474) );
  NAND3X1TF U924 ( .A(N893), .B(N198), .C(N197), .Y(N674) );
  NAND2X1TF U925 ( .A(N88), .B(C152_DATA4_8), .Y(N197) );
  OAI2BB1X1TF U926 ( .A0N(N88), .A1N(C152_DATA4_10), .B0(N199), .Y(N672) );
  AOI2BB1X1TF U927 ( .A0N(N511), .A1N(N484), .B0(N514), .Y(N485) );
  OR3X1TF U928 ( .A(N906), .B(N74), .C(N896), .Y(N190) );
  NAND3X1TF U929 ( .A(SIGN_Y), .B(N74), .C(N895), .Y(N823) );
  NAND2X1TF U930 ( .A(N892), .B(N859), .Y(N856) );
  CMPR32X2TF U931 ( .A(X_IN[1]), .B(DIVISION_HEAD[5]), .C(INTADD_0_CI), .CO(
        INTADD_0_N7), .S(\INTADD_0_SUM[0] ) );
  AOI2BB2X1TF U932 ( .B0(N205), .B1(DIVISION_REMA[0]), .A0N(N153), .A1N(N52), 
        .Y(N208) );
  OAI222X1TF U933 ( .A0(N54), .A1(N44), .B0(N52), .B1(N40), .C0(N227), .C1(
        N136), .Y(FOUT[10]) );
  OAI222X1TF U934 ( .A0(N227), .A1(N39), .B0(N52), .B1(N43), .C0(N133), .C1(
        N54), .Y(FOUT[9]) );
  NAND2X1TF U935 ( .A(N147), .B(N120), .Y(N370) );
  NAND3X1TF U936 ( .A(N545), .B(N387), .C(N634), .Y(N647) );
  AOI222XLTF U937 ( .A0(STEP[2]), .A1(N149), .B0(N121), .B1(N120), .C0(N134), 
        .C1(N122), .Y(N246) );
  NAND2X1TF U938 ( .A(N137), .B(N160), .Y(N616) );
  NAND2X1TF U939 ( .A(N565), .B(N956), .Y(N942) );
  NAND2X1TF U940 ( .A(N965), .B(N378), .Y(N573) );
  NOR2BX1TF U941 ( .AN(N573), .B(N605), .Y(N570) );
  NAND2X1TF U942 ( .A(PRE_WORK), .B(N351), .Y(N951) );
  NAND2X1TF U943 ( .A(N204), .B(N957), .Y(N363) );
  XNOR2X1TF U944 ( .A(OPER_A[12]), .B(N340), .Y(N341) );
  NAND3X1TF U945 ( .A(N605), .B(N602), .C(N141), .Y(N600) );
  NAND3X1TF U946 ( .A(N566), .B(POST_WORK), .C(N602), .Y(N373) );
  NAND3BX1TF U947 ( .AN(N363), .B(N950), .C(N965), .Y(N598) );
  NAND3X1TF U948 ( .A(N609), .B(N364), .C(N598), .Y(N945) );
  NAND2X1TF U949 ( .A(N75), .B(N395), .Y(N382) );
  NAND3X1TF U950 ( .A(N385), .B(N122), .C(DP_OP_333_124_4748_N57), .Y(N638) );
  NAND3BX1TF U951 ( .AN(N382), .B(N774), .C(N638), .Y(N366) );
  NOR2BX1TF U952 ( .AN(N634), .B(N946), .Y(N542) );
  NAND3X1TF U953 ( .A(N542), .B(N377), .C(N376), .Y(N381) );
  NAND2X1TF U954 ( .A(N798), .B(SUM_AB[8]), .Y(N425) );
  NAND4X1TF U955 ( .A(N428), .B(N427), .C(N426), .D(N425), .Y(N429) );
  NAND4X1TF U956 ( .A(N439), .B(N438), .C(N437), .D(N436), .Y(N440) );
  NAND4X1TF U957 ( .A(N449), .B(N448), .C(N447), .D(N446), .Y(N450) );
  AOI2BB2X1TF U958 ( .B0(X_IN[9]), .B1(N479), .A0N(N479), .A1N(X_IN[9]), .Y(
        N484) );
  NAND3X1TF U959 ( .A(N509), .B(N39), .C(N484), .Y(N480) );
  AOI2BB2X1TF U960 ( .B0(N488), .B1(N503), .A0N(N503), .A1N(N488), .Y(N495) );
  AOI2BB1X1TF U961 ( .A0N(N511), .A1N(N495), .B0(N514), .Y(N496) );
  AOI2BB2X1TF U962 ( .B0(X_IN[11]), .B1(N498), .A0N(N498), .A1N(X_IN[11]), .Y(
        N510) );
  OAI2BB2XLTF U963 ( .B0(N503), .B1(N608), .A0N(XTEMP[12]), .A1N(N502), .Y(
        N504) );
  AOI2BB1X1TF U964 ( .A0N(N511), .A1N(N510), .B0(N514), .Y(N512) );
  AOI2BB1X1TF U965 ( .A0N(DIVISION_REMA[2]), .A1N(N518), .B0(DIVISION_HEAD[6]), 
        .Y(N516) );
  OA21XLTF U966 ( .A0(N130), .A1(DIVISION_REMA[4]), .B0(N520), .Y(N522) );
  OA21XLTF U967 ( .A0(N132), .A1(DIVISION_REMA[6]), .B0(N524), .Y(N526) );
  OA21XLTF U968 ( .A0(XTEMP[12]), .A1(N535), .B0(N40), .Y(N534) );
  NAND4X1TF U969 ( .A(N545), .B(N544), .C(N638), .D(N543), .Y(N556) );
  NAND3X1TF U970 ( .A(N551), .B(N550), .C(N549), .Y(N552) );
  NAND3X1TF U971 ( .A(N754), .B(N559), .C(N558), .Y(N560) );
  NAND3X1TF U972 ( .A(N566), .B(N602), .C(N821), .Y(N572) );
  NAND4X1TF U973 ( .A(N568), .B(N567), .C(N639), .D(N572), .Y(N569) );
  NAND2X1TF U974 ( .A(N159), .B(N138), .Y(N590) );
  NOR4XLTF U975 ( .A(\RSHT_BITS[3] ), .B(N90), .C(N614), .D(N590), .Y(N571) );
  NAND2X1TF U976 ( .A(N579), .B(N589), .Y(N586) );
  NAND2X1TF U977 ( .A(N92), .B(N91), .Y(N588) );
  AOI2BB2X1TF U978 ( .B0(N596), .B1(N138), .A0N(N590), .A1N(N592), .Y(N584) );
  NAND4X1TF U979 ( .A(N611), .B(N610), .C(N609), .D(N608), .Y(N612) );
  NAND4X1TF U980 ( .A(N47), .B(N634), .C(N633), .D(N632), .Y(N635) );
  NAND4X1TF U981 ( .A(N640), .B(N639), .C(N638), .D(N643), .Y(N697) );
  NAND3X1TF U982 ( .A(N754), .B(N651), .C(N650), .Y(N652) );
  AO22X1TF U983 ( .A0(DIVISION_REMA[4]), .A1(N80), .B0(N172), .B1(N788), .Y(
        N742) );
  NAND4X1TF U984 ( .A(N792), .B(N791), .C(N790), .D(N789), .Y(N793) );
  OAI221XLTF U985 ( .A0(\INDEX[2] ), .A1(N90), .B0(N124), .B1(\RSHT_BITS[3] ), 
        .C0(N816), .Y(N817) );
  OAI221XLTF U986 ( .A0(N129), .A1(N159), .B0(N137), .B1(N92), .C0(N818), .Y(
        N832) );
  NAND2X1TF U987 ( .A(N831), .B(N965), .Y(N860) );
  NAND3X1TF U988 ( .A(SIGN_Y), .B(N74), .C(N206), .Y(N835) );
  OAI2BB1X1TF U989 ( .A0N(N958), .A1N(N832), .B0(N831), .Y(N916) );
  NAND3X1TF U990 ( .A(N74), .B(N157), .C(N45), .Y(N973) );
  NAND3BX1TF U991 ( .AN(OPER_A[7]), .B(N928), .C(N879), .Y(N880) );
  NAND3X1TF U992 ( .A(N905), .B(N904), .C(N903), .Y(N673) );
  NAND2X1TF U993 ( .A(N978), .B(N977), .Y(N668) );
  NAND2X1TF U994 ( .A(N981), .B(N980), .Y(N667) );
  NAND2X1TF U995 ( .A(SUM_AB[3]), .B(N49), .Y(N982) );
  NAND2X1TF U996 ( .A(N987), .B(N986), .Y(N665) );
  NAND2X1TF U997 ( .A(SUM_AB[5]), .B(N171), .Y(N988) );
  NAND2X1TF U998 ( .A(N993), .B(N992), .Y(N663) );
  NAND2X1TF U999 ( .A(SUM_AB[7]), .B(N171), .Y(N994) );
  NAND2X1TF U1000 ( .A(N999), .B(N998), .Y(N661) );
  NAND2X1TF U1001 ( .A(SUM_AB[9]), .B(N171), .Y(N1000) );
  NAND2X1TF U1002 ( .A(N1005), .B(N1004), .Y(N659) );
  NAND2X1TF U1003 ( .A(SUM_AB[11]), .B(N171), .Y(N1006) );
endmodule


module SERIAL_CPU_8BIT_VG ( CLK, ENABLE, RST_N, START, I_DATAIN, D_DATAIN, 
        IS_I_ADDR, NXT, I_ADDR, D_ADDR, D_WE, D_DATAOUT, IO_STATUS, IO_CONTROL, 
        IO_DATAINA, IO_DATAINB, IO_DATAOUTA, IO_DATAOUTB, IO_OFFSET );
  input [7:0] I_DATAIN;
  input [7:0] D_DATAIN;
  output [1:0] NXT;
  output [8:0] I_ADDR;
  output [8:0] D_ADDR;
  output [7:0] D_DATAOUT;
  input [15:0] IO_STATUS;
  output [15:0] IO_CONTROL;
  input [15:0] IO_DATAINA;
  input [15:0] IO_DATAINB;
  output [15:0] IO_DATAOUTA;
  output [15:0] IO_DATAOUTB;
  output [15:0] IO_OFFSET;
  input CLK, ENABLE, RST_N, START;
  output IS_I_ADDR, D_WE;
  wire   N163, N164, N165, CF_BUF, N467, N468, N469, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N501,
         N502, N503, N504, N505, N506, N507, N508, N509, N510, N511, N512,
         N513, N514, N515, N516, N517, N585, N586, ZF, NF, CF, N403, N411,
         N412, N413, N414, N415, N417, N418, N419, N425, N427, N446, N448,
         N450, N451, N452, N453, N454, N455, N456, N457, N458, N459, N460,
         N463, N464, N465, N466, N4730, N4750, N4770, N4780, N4800, N4810,
         N4830, N484, N486, N5110, N5120, N5130, N5140, N5150, N5160, N5170,
         N518, N519, N520, N521, N522, N524, N526, N528, N530, N532, N534,
         N536, N538, N573, N575, N577, N579, N581, N583, N5850, N587, N589,
         N593, N594, N597, N598, N601, N602, N605, N606, N609, N610, N613,
         N614, N617, N618, N621, N622, N625, N626, N629, N633, N634, N637,
         N638, N641, N642, N645, N651, N654, N655, N656, N657, N658, N659,
         N660, N661, N679, N693, N695, N696, N697, N720, N721, N722, N723,
         N724, N725, N726, N727, N728, N729, N730, N731, N732, N733, N734,
         N735, N738, N739, N740, N741, N742, N743, N744, N745, N746, N747,
         N748, N749, N750, N751, N752, N753, N754, N755, N756, N757, N758,
         N759, N760, N761, N762, N763, N764, N765, N766, N767, N768, N769,
         N770, N771, N772, N773, N774, N775, N776, N777, N778, N779, N780,
         N781, N782, N783, N784, N785, N786, N787, N788, N789, N790, N791,
         N792, N793, N794, N795, N796, N797, N798, N799, N800, N801, N802,
         N803, N804, N805, N806, N807, N808, N809, N810, N811, N812, N813,
         N814, N815, N816, N817, N1050, N1051, N1052, N1053, N1054, N1055,
         N1056, N1057, N1058, N1059, N1060, N1061, N1062, N1063, N1064, N1065,
         N1066, N1067, N1068, N1069, N1070, N1071, N1072, N1073, N1074, N1075,
         N1076, N1077, N1078, N1079, N1080, N1081, N1082, N1083, N1084, N1085,
         N1086, N1087, N1088, N1089, N1090, N1091, N1092, N1093, N1094, N1095,
         N1096, N1097, N1098, N1099, N1100, N1101, N1102, N1103, N1104, N1105,
         N1106, N1107, N1108, N1109, N1110, N1111, N1112, N1113, N1114, N1115,
         N1116, N1117, N1118, N1119, N1120, N1121, N1122, N1123, N1124, N1125,
         N1126, N1127, N1128, N1129, N1130, N1131, ADD_X_276_3_N22,
         ADD_X_276_3_N21, ADD_X_276_3_N20, ADD_X_276_3_N19, ADD_X_276_3_N18,
         ADD_X_276_3_N17, ADD_X_276_3_N16, ADD_X_276_3_N15, ADD_X_276_3_N14,
         ADD_X_276_3_N13, ADD_X_276_3_N12, ADD_X_276_3_N11, ADD_X_276_3_N10,
         ADD_X_276_3_N9, ADD_X_276_3_N8, ADD_X_276_3_N7, ADD_X_276_3_N6,
         ADD_X_276_3_N5, ADD_X_276_3_N4, ADD_X_276_3_N3, ADD_X_276_3_N2,
         \SUB_X_276_4_B[0] , SUB_X_276_4_N16, SUB_X_276_4_N15, SUB_X_276_4_N14,
         SUB_X_276_4_N13, SUB_X_276_4_N12, SUB_X_276_4_N11, SUB_X_276_4_N10,
         SUB_X_276_4_N9, SUB_X_276_4_N8, SUB_X_276_4_N7, SUB_X_276_4_N6,
         SUB_X_276_4_N5, SUB_X_276_4_N4, SUB_X_276_4_N3, SUB_X_276_4_N2,
         SUB_X_276_4_N1, N1, N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12,
         N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23, N24, N25, N26,
         N27, N28, N29, N30, N31, N32, N33, N34, N35, N36, N37, N38, N39, N40,
         N41, N42, N43, N44, N45, N46, N47, N48, N49, N50, N51, N52, N53, N54,
         N55, N56, N57, N58, N59, N60, N97, N159, N160, N161, N162, N1630,
         N1640, N1650, N166, N167, N168, N169, N170, N171, N172, N173, N174,
         N175, N176, N177, N178, N179, N180, N181, N182, N183, N184, N186,
         N187, N188, N189, N190, N191, N192, N193, N194, N195, N196, N197,
         N198, N199, N200, N201, N202, N203, N204, N205, N206, N207, N208,
         N209, N210, N211, N212, N213, N214, N215, N216, N217, N218, N219,
         N220, N221, N222, N223, N259, N260, N261, N262, N263, N264, N265,
         N266, N267, N268, N269, N270, N271, N272, N273, N274, N275, N276,
         N277, N278, N279, N280, N281, N282, N283, N284, N285, N286, N287,
         N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298,
         N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N309,
         N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320,
         N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331,
         N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342,
         N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353,
         N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, N364,
         N365, N366, N367, N368, N369, N370, N371, N372, N373, N374, N375,
         N376, N377, N378, N379, N380, N381, N382, N383, N384, N385, N386,
         N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397,
         N398, N399, N400, N401, N402, N404, N405, N406, N407, N408, N409,
         N410, N416, N420, N421, N422, N423, N424, N426, N428, N429, N430,
         N431, N432, N433, N434, N435, N436, N437, N438, N439, N440, N441,
         N442, N443, N444, N445, N447, N449, N461, N462, N4670, N4680, N4690,
         N4700, N4710, N4720, N4740, N4760, N4790, N4820, N485, N487, N488,
         N489, N490, N491, N492, N493, N494, N495, N496, N497, N498, N499,
         N500, N5010, N5020, N5030, N5040, N5050, N5060, N5070, N5080, N5090,
         N5100, N523, N525, N527, N529, N531, N533, N535, N537, N539, N540,
         N541, N542, N543, N544, N545, N546, N547, N548, N549, N550, N551,
         N552, N553, N554, N555, N556, N557, N558, N559, N560, N561, N562,
         N563, N564, N565, N566, N567, N568, N569, N570, N571, N572, N574,
         N576, N578, N580, N582, N584, N5860, N588, N590, N591, N592, N595,
         N596, N599, N600, N603, N604, N607, N608, N611, N612, N615, N616,
         N619, N620, N623, N624, N627, N628, N630, N631, N632, N635, N636,
         N639, N640, N643, N644, N646, N647, N648, N650, N652, N653, N662,
         N663, N664, N665, N666, N667, N668, N669, N670, N671, N672, N673,
         N674, N675, N676, N677, N678, N680, N681, N682, N683, N684, N685,
         N686, N687, N688, N689, N690, N691, N692, N694, N698, N699, N700,
         N701, N702, N703, N704, N705, N706, N707, N708, N709, N710, N711,
         N712, N713, N714, N715, N716, N717, N718, N719, N736, N737, N818,
         N819, N820, N821, N822, N823, N824, N825, N826, N827, N828, N829,
         N830, N831, N832, N833, N834, N835, N836, N837, N838, N839, N840,
         N841, N842, N843, N844, N845, N846, N847, N848, N849, N850, N851,
         N852, N853, N854, N855, N856, N857, N858, N859, N860, N861, N862,
         N863, N864, N865, N866, N867, N868, N869, N870, N871, N872, N873,
         N874, N875, N876, N877, N878, N879, N880, N881, N882, N883, N884,
         N885, N886, N887, N888, N889, N890, N891, N892, N893, N894, N895,
         N896, N897, N898, N899, N900, N901, N902, N903, N904, N905, N906,
         N907, N908, N909, N910, N911, N912, N913, N914, N915, N916, N917,
         N918, N919, N920, N921, N922, N923, N924, N925, N926, N927, N928,
         N929, N930, N931, N932, N933, N934, N935, N936, N937, N938, N939,
         N940, N941, N942, N943, N944, N945, N946, N947, N948, N949, N950,
         N951, N952, N953, N954, N955, N956, N957, N958, N959, N960, N961,
         N962, N963, N964, N965, N966, N967, N968, N969, N970, N971, N972,
         N973, N974, N975, N976, N977, N978, N979, N980, N981, N982, N983,
         N984, N985, N986, N987, N988, N989, N990, N991, N992, N993, N994,
         N995, N996, N997, N998, N999, N1000, N1001, N1002, N1003, N1004,
         N1005, N1006, N1007, N1008, N1009, N1010, N1011, N1012, N1013, N1014,
         N1015, N1016, N1017, N1018, N1019, N1020, N1021, N1022, N1023, N1024,
         N1025, N1026, N1027, N1028, N1029, N1030, N1031, N1032, N1033, N1034,
         N1035, N1036, N1037, N1038, N1039, N1040, N1041, N1042, N1043, N1044,
         N1045, N1046, N1047, N1048, N1049, N1132, N1133, N1134, N1135, N1136,
         N1137, N1138, N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1146,
         N1147, N1148, N1149, N1150, N1151, N1152, N1153, N1154, N1155, N1156,
         N1157, N1158, N1159, N1160, N1161, N1162, N1163, N1164, N1165, N1166,
         N1167, N1168, N1169, N1170, N1171, N1172, N1173, N1174, N1175, N1176,
         N1177, N1178, N1179, N1180, N1181, N1182, N1183, N1184, N1185, N1186,
         N1187, N1188, N1189, N1190, N1191, N1192, N1193, N1194, N1195, N1196,
         N1197, N1198, N1199, N1200, N1201, N1202, N1203, N1204, N1205, N1206,
         N1207, N1208, N1209, N1210, N1211, N1212, N1213, N1214, N1215, N1216,
         N1217, N1218, N1219, N1220, N1221, N1222, N1223, N1224, N1225, N1226,
         N1227, N1228, N1229, N1230, N1231, N1232, N1233, N1234, N1235, N1236,
         N1237, N1238;
  wire   [3:1] STATE;
  wire   [4:2] CODE_TYPE;
  wire   [2:0] OPER3_R3;
  wire   [2:0] NEXT_STATE;
  wire   [15:0] REG_A;
  wire   [15:0] REG_B;
  wire   [15:14] REG_C;

  DFFNSRX4TF \gr_reg[3][0]  ( .D(N1065), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_DATAOUTB[0]), .QN(N769) );
  DFFNSRX4TF \gr_reg[3][1]  ( .D(N1064), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_DATAOUTB[1]), .QN(N768) );
  DFFNSRX4TF \gr_reg[3][2]  ( .D(N1063), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_DATAOUTB[2]), .QN(N767) );
  AFCSIHCONX2TF \add_x_276_3/U17  ( .A(REG_B[2]), .B(REG_A[2]), .CS(
        ADD_X_276_3_N21), .S(N469), .CO0N(ADD_X_276_3_N20), .CO1N(
        ADD_X_276_3_N19) );
  AFCSHCINX2TF \add_x_276_3/U16  ( .CI1N(ADD_X_276_3_N19), .B(REG_B[3]), .A(
        REG_A[3]), .CI0N(ADD_X_276_3_N20), .CS(ADD_X_276_3_N21), .CO1(
        ADD_X_276_3_N17), .CO0(ADD_X_276_3_N18), .S(N470) );
  AFCSIHCONX2TF \add_x_276_3/U14  ( .A(REG_A[4]), .B(REG_B[4]), .CS(
        ADD_X_276_3_N16), .S(N471), .CO0N(ADD_X_276_3_N15), .CO1N(
        ADD_X_276_3_N14) );
  AFCSHCINX2TF \add_x_276_3/U13  ( .CI1N(ADD_X_276_3_N14), .B(REG_A[5]), .A(
        REG_B[5]), .CI0N(ADD_X_276_3_N15), .CS(ADD_X_276_3_N16), .CO1(
        ADD_X_276_3_N12), .CO0(ADD_X_276_3_N13), .S(N472) );
  CMPR32X2TF \add_x_276_3/U11  ( .A(REG_A[6]), .B(REG_B[6]), .C(
        ADD_X_276_3_N11), .CO(ADD_X_276_3_N10), .S(N473) );
  CMPR32X2TF \add_x_276_3/U10  ( .A(REG_A[7]), .B(REG_B[7]), .C(
        ADD_X_276_3_N10), .CO(ADD_X_276_3_N9), .S(N474) );
  CMPR32X2TF \add_x_276_3/U9  ( .A(REG_A[8]), .B(REG_B[8]), .C(ADD_X_276_3_N9), 
        .CO(ADD_X_276_3_N8), .S(N475) );
  CMPR32X2TF \add_x_276_3/U8  ( .A(REG_A[9]), .B(REG_B[9]), .C(ADD_X_276_3_N8), 
        .CO(ADD_X_276_3_N7), .S(N476) );
  CMPR32X2TF \add_x_276_3/U7  ( .A(REG_A[10]), .B(REG_B[10]), .C(
        ADD_X_276_3_N7), .CO(ADD_X_276_3_N6), .S(N477) );
  CMPR32X2TF \add_x_276_3/U6  ( .A(REG_A[11]), .B(REG_B[11]), .C(
        ADD_X_276_3_N6), .CO(ADD_X_276_3_N5), .S(N478) );
  CMPR32X2TF \add_x_276_3/U5  ( .A(REG_A[12]), .B(REG_B[12]), .C(
        ADD_X_276_3_N5), .CO(ADD_X_276_3_N4), .S(N479) );
  CMPR32X2TF \add_x_276_3/U4  ( .A(REG_A[13]), .B(REG_B[13]), .C(
        ADD_X_276_3_N4), .CO(ADD_X_276_3_N3), .S(N480) );
  CMPR32X2TF \add_x_276_3/U3  ( .A(REG_A[14]), .B(REG_B[14]), .C(
        ADD_X_276_3_N3), .CO(ADD_X_276_3_N2), .S(N481) );
  DFFNSRX2TF nf_reg ( .D(N448), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(NF), .QN(
        N294) );
  DFFNSRX2TF \pc_reg[7]  ( .D(N655), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        I_ADDR[8]), .QN(N293) );
  DFFNSRX2TF \pc_reg[0]  ( .D(N654), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        I_ADDR[1]), .QN(N292) );
  DFFNSRX2TF \state_reg[0]  ( .D(NEXT_STATE[0]), .CKN(CLK), .SN(1'b1), .RN(
        RST_N), .Q(N291), .QN(N679) );
  DFFNSRX2TF zf_reg ( .D(N450), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(ZF), .QN(
        N290) );
  DFFNSRX2TF \gr_reg[3][12]  ( .D(N1101), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .Q(IO_DATAOUTB[12]), .QN(N757) );
  DFFNSRX2TF \gr_reg[4][0]  ( .D(N1057), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_OFFSET[0]), .QN(N753) );
  DFFNSRX2TF \gr_reg[4][1]  ( .D(N1056), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_OFFSET[1]), .QN(N752) );
  DFFNSRX2TF \gr_reg[4][2]  ( .D(N1055), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_OFFSET[2]), .QN(N751) );
  DFFNSRX2TF \gr_reg[4][3]  ( .D(N1054), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_OFFSET[3]), .QN(N750) );
  DFFNSRX2TF \gr_reg[4][5]  ( .D(N1052), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_OFFSET[5]), .QN(N748) );
  DFFNSRX2TF \gr_reg[4][7]  ( .D(N1050), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_OFFSET[7]), .QN(N746) );
  DFFNSRX2TF \gr_reg[2][2]  ( .D(N1071), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_DATAOUTA[2]), .QN(N783) );
  DFFNSRX2TF \gr_reg[2][5]  ( .D(N1068), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_DATAOUTA[5]), .QN(N780) );
  DFFNSRX2TF \gr_reg[2][7]  ( .D(N1066), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_DATAOUTA[7]), .QN(N778) );
  DFFNSRX2TF \gr_reg[3][5]  ( .D(N1060), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_DATAOUTB[5]), .QN(N764) );
  DFFNSRX2TF \gr_reg[3][14]  ( .D(N1099), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .Q(N286), .QN(N755) );
  DFFNSRX2TF \gr_reg[3][13]  ( .D(N1100), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .Q(N285), .QN(N756) );
  DFFNSRX2TF \gr_reg[3][4]  ( .D(N1061), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_DATAOUTB[4]), .QN(N765) );
  DFFNSRX2TF \gr_reg[3][6]  ( .D(N1059), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_DATAOUTB[6]), .QN(N763) );
  DFFNSRX2TF \gr_reg[3][8]  ( .D(N1105), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_DATAOUTB[8]), .QN(N761) );
  DFFNSRX2TF \gr_reg[3][10]  ( .D(N1103), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .Q(IO_DATAOUTB[10]), .QN(N759) );
  DFFNSRX2TF \gr_reg[3][11]  ( .D(N1102), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .Q(IO_DATAOUTB[11]), .QN(N758) );
  DFFNSRX2TF \gr_reg[3][15]  ( .D(N1098), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .Q(N284), .QN(N754) );
  DFFNSRX2TF \id_ir_reg[5]  ( .D(N534), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        N281), .QN(N413) );
  DFFNSRX2TF \id_ir_reg[14]  ( .D(N577), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        CODE_TYPE[3]), .QN(N264) );
  DFFNSRX2TF \id_ir_reg[9]  ( .D(N587), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        N275), .QN(N696) );
  DFFNSRX2TF \state_reg[1]  ( .D(NEXT_STATE[1]), .CKN(CLK), .SN(1'b1), .RN(
        RST_N), .Q(STATE[1]), .QN(N270) );
  DFFNSRX2TF \gr_reg[2][1]  ( .D(N1072), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_DATAOUTA[1]), .QN(N784) );
  DFFNSRX2TF \gr_reg[2][3]  ( .D(N1070), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_DATAOUTA[3]), .QN(N782) );
  DFFNSRX2TF \gr_reg[3][7]  ( .D(N1058), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_DATAOUTB[7]), .QN(N762) );
  DFFNSRX2TF \id_ir_reg[2]  ( .D(N528), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        OPER3_R3[2]), .QN(N269) );
  DFFNSRX2TF \state_reg[2]  ( .D(NEXT_STATE[2]), .CKN(CLK), .SN(1'b1), .RN(
        RST_N), .Q(STATE[2]), .QN(N268) );
  DFFNSRX2TF \id_ir_reg[10]  ( .D(N5850), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .Q(N265), .QN(N695) );
  DFFNSRX2TF \id_ir_reg[15]  ( .D(N575), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        CODE_TYPE[4]), .QN(N263) );
  DFFNSRX2TF \id_ir_reg[1]  ( .D(N526), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        OPER3_R3[1]), .QN(N261) );
  DFFNSRX2TF \id_ir_reg[8]  ( .D(N589), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        N260), .QN(N697) );
  DFFNSRX2TF \id_ir_reg[0]  ( .D(N524), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        OPER3_R3[0]), .QN(N259) );
  TLATXLTF cf_buf_reg ( .G(N585), .D(N586), .Q(CF_BUF) );
  TLATXLTF \nxt_reg[0]  ( .G(N163), .D(N164), .Q(NXT[0]) );
  TLATXLTF \nxt_reg[1]  ( .G(N163), .D(N165), .Q(NXT[1]) );
  DFFRX2TF \smdr_reg[0]  ( .D(N486), .CK(CLK), .RN(RST_N), .QN(N735) );
  DFFRX2TF \smdr_reg[1]  ( .D(N4830), .CK(CLK), .RN(RST_N), .QN(N734) );
  DFFRX2TF \smdr_reg[2]  ( .D(N4800), .CK(CLK), .RN(RST_N), .QN(N733) );
  DFFRX2TF \smdr_reg[3]  ( .D(N4770), .CK(CLK), .RN(RST_N), .QN(N732) );
  DFFRX2TF \smdr_reg[4]  ( .D(N4750), .CK(CLK), .RN(RST_N), .QN(N731) );
  DFFRX2TF \smdr_reg[6]  ( .D(N4730), .CK(CLK), .RN(RST_N), .QN(N729) );
  DFFRX2TF \smdr_reg[5]  ( .D(N466), .CK(CLK), .RN(RST_N), .QN(N730) );
  DFFRX2TF \smdr_reg[7]  ( .D(N460), .CK(CLK), .RN(RST_N), .QN(N728) );
  DFFRX2TF \smdr_reg[8]  ( .D(N522), .CK(CLK), .RN(RST_N), .QN(N727) );
  DFFRX2TF \smdr_reg[9]  ( .D(N521), .CK(CLK), .RN(RST_N), .QN(N726) );
  DFFRX2TF \smdr_reg[10]  ( .D(N520), .CK(CLK), .RN(RST_N), .QN(N725) );
  DFFRX2TF \smdr_reg[11]  ( .D(N519), .CK(CLK), .RN(RST_N), .QN(N724) );
  DFFRX2TF \smdr_reg[12]  ( .D(N518), .CK(CLK), .RN(RST_N), .QN(N723) );
  DFFRX2TF \smdr_reg[13]  ( .D(N5170), .CK(CLK), .RN(RST_N), .QN(N722) );
  DFFRX2TF \smdr_reg[14]  ( .D(N5160), .CK(CLK), .RN(RST_N), .QN(N721) );
  DFFRX2TF \smdr_reg[15]  ( .D(N5150), .CK(CLK), .RN(RST_N), .QN(N720) );
  DFFNSRX2TF \reg_C_reg[14]  ( .D(N637), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_C[14]) );
  DFFNSRX2TF \reg_C_reg[15]  ( .D(N645), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        REG_C[15]) );
  DFFNSRX2TF cf_reg ( .D(N446), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(CF) );
  DFFNSRX2TF \gr_reg[4][8]  ( .D(N1097), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_OFFSET[8]), .QN(N745) );
  DFFNSRX2TF \gr_reg[4][9]  ( .D(N1096), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_OFFSET[9]), .QN(N744) );
  DFFNSRX2TF \pc_reg[6]  ( .D(N661), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        I_ADDR[7]) );
  DFFNSRX2TF \pc_reg[4]  ( .D(N659), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        I_ADDR[5]) );
  DFFNSRX2TF \reg_C_reg[1]  ( .D(N633), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        D_ADDR[2]) );
  DFFNSRX2TF \reg_C_reg[3]  ( .D(N617), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        D_ADDR[4]) );
  DFFNSRX2TF \reg_C_reg[4]  ( .D(N609), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        D_ADDR[5]) );
  DFFNSRX2TF \reg_C_reg[6]  ( .D(N605), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        D_ADDR[7]) );
  DFFNSRX2TF \reg_C_reg[2]  ( .D(N597), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        D_ADDR[3]) );
  DFFNSRX2TF \reg_C_reg[7]  ( .D(N593), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        D_ADDR[8]) );
  DFFNSRX2TF \reg_C_reg[5]  ( .D(N463), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        D_ADDR[6]) );
  DFFNSRX2TF \pc_reg[2]  ( .D(N657), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        I_ADDR[3]) );
  DFFNSRX2TF \pc_reg[5]  ( .D(N660), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        I_ADDR[6]) );
  DFFNSRX2TF \pc_reg[3]  ( .D(N658), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        I_ADDR[4]) );
  DFFNSRX2TF \pc_reg[1]  ( .D(N656), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        I_ADDR[2]) );
  DFFNSRX2TF \gr_reg[4][4]  ( .D(N1053), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_OFFSET[4]), .QN(N749) );
  DFFNSRX2TF \gr_reg[4][6]  ( .D(N1051), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_OFFSET[6]), .QN(N747) );
  DFFNSRX2TF \gr_reg[1][0]  ( .D(N1081), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_CONTROL[0]), .QN(N801) );
  DFFNSRX2TF \gr_reg[2][11]  ( .D(N1110), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .Q(IO_DATAOUTA[11]), .QN(N774) );
  DFFNSRX2TF \gr_reg[1][1]  ( .D(N1080), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_CONTROL[1]), .QN(N800) );
  DFFNSRX2TF \gr_reg[2][12]  ( .D(N1109), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .Q(IO_DATAOUTA[12]), .QN(N773) );
  DFFNSRX2TF \gr_reg[2][10]  ( .D(N1111), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .Q(IO_DATAOUTA[10]), .QN(N775) );
  DFFRX2TF \reg_B_reg[0]  ( .D(N638), .CK(CLK), .RN(RST_N), .Q(REG_B[0]), .QN(
        N54) );
  DFFRX2TF \reg_B_reg[2]  ( .D(N594), .CK(CLK), .RN(RST_N), .Q(REG_B[2]), .QN(
        N57) );
  DFFNSRX2TF \gr_reg[1][5]  ( .D(N1076), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_CONTROL[5]), .QN(N796) );
  DFFNSRX2TF \gr_reg[2][4]  ( .D(N1069), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_DATAOUTA[4]), .QN(N781) );
  DFFNSRX2TF \gr_reg[1][2]  ( .D(N1079), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_CONTROL[2]), .QN(N799) );
  DFFNSRX2TF \gr_reg[1][4]  ( .D(N1077), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_CONTROL[4]), .QN(N797) );
  DFFNSRX2TF \gr_reg[1][3]  ( .D(N1078), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_CONTROL[3]), .QN(N798) );
  DFFNSRX2TF \gr_reg[3][9]  ( .D(N1104), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_DATAOUTB[9]), .QN(N760) );
  DFFRX2TF \reg_A_reg[1]  ( .D(N484), .CK(CLK), .RN(RST_N), .Q(REG_A[1]), .QN(
        N59) );
  DFFNSRX2TF \id_ir_reg[13]  ( .D(N579), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        CODE_TYPE[2]), .QN(N55) );
  DFFNSRX2TF \gr_reg[2][8]  ( .D(N1113), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_DATAOUTA[8]), .QN(N777) );
  DFFNSRX2TF \gr_reg[3][3]  ( .D(N1062), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_DATAOUTB[3]), .QN(N766) );
  DFFNSRX2TF \gr_reg[2][9]  ( .D(N1112), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_DATAOUTA[9]), .QN(N776) );
  DFFNSRX2TF \id_ir_reg[12]  ( .D(N581), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        N289), .QN(N693) );
  ADDHXLTF \add_x_276_3/U19  ( .A(\SUB_X_276_4_B[0] ), .B(REG_A[0]), .CO(
        ADD_X_276_3_N22), .S(N467) );
  CMPR32X2TF \add_x_276_3/U2  ( .A(REG_A[15]), .B(REG_B[15]), .C(
        ADD_X_276_3_N2), .CO(N483), .S(N482) );
  CMPR32X2TF \add_x_276_3/U18  ( .A(REG_A[1]), .B(REG_B[1]), .C(
        ADD_X_276_3_N22), .CO(ADD_X_276_3_N21), .S(N468) );
  CLKMX2X2TF \add_x_276_3/U12  ( .A(ADD_X_276_3_N13), .B(ADD_X_276_3_N12), 
        .S0(ADD_X_276_3_N16), .Y(ADD_X_276_3_N11) );
  DFFNSRX4TF \gr_reg[2][0]  ( .D(N1073), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_DATAOUTA[0]), .QN(N785) );
  CMPR32X2TF \sub_x_276_4/U10  ( .A(N215), .B(REG_A[7]), .C(SUB_X_276_4_N10), 
        .CO(SUB_X_276_4_N9), .S(N508) );
  CMPR32X2TF \sub_x_276_4/U14  ( .A(N60), .B(REG_A[3]), .C(SUB_X_276_4_N14), 
        .CO(SUB_X_276_4_N13), .S(N504) );
  CMPR32X2TF \sub_x_276_4/U15  ( .A(N57), .B(REG_A[2]), .C(SUB_X_276_4_N15), 
        .CO(SUB_X_276_4_N14), .S(N503) );
  CMPR32X2TF \sub_x_276_4/U8  ( .A(N217), .B(REG_A[9]), .C(SUB_X_276_4_N8), 
        .CO(SUB_X_276_4_N7), .S(N510) );
  CMPR32X2TF \sub_x_276_4/U6  ( .A(N219), .B(REG_A[11]), .C(SUB_X_276_4_N6), 
        .CO(SUB_X_276_4_N5), .S(N512) );
  CMPR32X2TF \sub_x_276_4/U12  ( .A(N213), .B(REG_A[5]), .C(SUB_X_276_4_N12), 
        .CO(SUB_X_276_4_N11), .S(N506) );
  CMPR32X2TF \sub_x_276_4/U11  ( .A(N214), .B(REG_A[6]), .C(SUB_X_276_4_N11), 
        .CO(SUB_X_276_4_N10), .S(N507) );
  CMPR32X2TF \sub_x_276_4/U13  ( .A(N212), .B(REG_A[4]), .C(SUB_X_276_4_N13), 
        .CO(SUB_X_276_4_N12), .S(N505) );
  CMPR32X2TF \sub_x_276_4/U9  ( .A(N216), .B(REG_A[8]), .C(SUB_X_276_4_N9), 
        .CO(SUB_X_276_4_N8), .S(N509) );
  CMPR32X2TF \sub_x_276_4/U7  ( .A(N218), .B(REG_A[10]), .C(SUB_X_276_4_N7), 
        .CO(SUB_X_276_4_N6), .S(N511) );
  CMPR32X2TF \sub_x_276_4/U5  ( .A(N220), .B(REG_A[12]), .C(SUB_X_276_4_N5), 
        .CO(SUB_X_276_4_N4), .S(N513) );
  CMPR32X2TF \sub_x_276_4/U3  ( .A(N222), .B(REG_A[14]), .C(SUB_X_276_4_N3), 
        .CO(SUB_X_276_4_N2), .S(N515) );
  CMPR32X2TF \sub_x_276_4/U4  ( .A(N221), .B(REG_A[13]), .C(SUB_X_276_4_N4), 
        .CO(SUB_X_276_4_N3), .S(N514) );
  DFFNSRX2TF \state_reg[3]  ( .D(N651), .CKN(CLK), .SN(RST_N), .RN(1'b1), .Q(
        N262), .QN(STATE[3]) );
  DFFNSRX2TF \gr_reg[2][6]  ( .D(N1067), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_DATAOUTA[6]), .QN(N779) );
  DFFNSRXLTF \reg_C_reg[8]  ( .D(N601), .CKN(CLK), .SN(1'b1), .RN(RST_N), .QN(
        N425) );
  DFFNSRXLTF \id_ir_reg[7]  ( .D(N538), .CKN(CLK), .SN(1'b1), .RN(RST_N), .QN(
        N403) );
  DFFNSRXLTF \id_ir_reg[3]  ( .D(N530), .CKN(CLK), .SN(1'b1), .RN(RST_N), .QN(
        N417) );
  DFFNSRXLTF \reg_C_reg[9]  ( .D(N613), .CKN(CLK), .SN(1'b1), .RN(RST_N), .QN(
        N419) );
  DFFNSRXLTF \reg_C_reg[10]  ( .D(N573), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N427) );
  DFFNSRXLTF \reg_C_reg[12]  ( .D(N621), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N418) );
  DFFNSRXLTF \reg_C_reg[11]  ( .D(N625), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N415) );
  DFFNSRXLTF \reg_C_reg[13]  ( .D(N629), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N414) );
  DFFNSRXLTF dw_reg ( .D(N1130), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(D_WE) );
  DFFNSRX2TF lowest_bit_reg ( .D(N1131), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        I_ADDR[0]), .QN(N288) );
  DFFNSRX2TF \reg_C_reg[0]  ( .D(N641), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        D_ADDR[1]) );
  DFFSX4TF \reg_A_reg[0]  ( .D(N97), .CK(CLK), .SN(RST_N), .Q(N1014), .QN(
        REG_A[0]) );
  DFFRX2TF \reg_B_reg[6]  ( .D(N456), .CK(CLK), .RN(RST_N), .Q(REG_B[6]), .QN(
        N214) );
  DFFRX2TF \reg_B_reg[5]  ( .D(N464), .CK(CLK), .RN(RST_N), .Q(REG_B[5]), .QN(
        N213) );
  DFFRX2TF \reg_B_reg[4]  ( .D(N455), .CK(CLK), .RN(RST_N), .Q(REG_B[4]), .QN(
        N212) );
  DFFRX2TF \reg_B_reg[3]  ( .D(N614), .CK(CLK), .RN(RST_N), .Q(REG_B[3]), .QN(
        N211) );
  DFFRX2TF \reg_B_reg[14]  ( .D(N451), .CK(CLK), .RN(RST_N), .Q(REG_B[14]), 
        .QN(N222) );
  DFFRX2TF \reg_B_reg[13]  ( .D(N452), .CK(CLK), .RN(RST_N), .Q(REG_B[13]), 
        .QN(N221) );
  DFFRX2TF \reg_B_reg[12]  ( .D(N453), .CK(CLK), .RN(RST_N), .Q(REG_B[12]), 
        .QN(N220) );
  DFFRX2TF \reg_A_reg[7]  ( .D(N459), .CK(CLK), .RN(RST_N), .Q(REG_A[7]), .QN(
        N272) );
  DFFRX2TF \reg_A_reg[5]  ( .D(N465), .CK(CLK), .RN(RST_N), .Q(REG_A[5]), .QN(
        N282) );
  DFFRX2TF \reg_A_reg[3]  ( .D(N4780), .CK(CLK), .RN(RST_N), .Q(REG_A[3]), 
        .QN(N273) );
  DFFRX2TF \reg_A_reg[2]  ( .D(N4810), .CK(CLK), .RN(RST_N), .Q(REG_A[2]), 
        .QN(N271) );
  DFFRX2TF \reg_B_reg[10]  ( .D(N5110), .CK(CLK), .RN(RST_N), .Q(REG_B[10]), 
        .QN(N218) );
  DFFRX2TF \reg_B_reg[7]  ( .D(N458), .CK(CLK), .RN(RST_N), .Q(REG_B[7]), .QN(
        N215) );
  DFFRX2TF \reg_B_reg[15]  ( .D(N642), .CK(CLK), .RN(RST_N), .Q(REG_B[15]), 
        .QN(N223) );
  DFFRX2TF \reg_B_reg[11]  ( .D(N622), .CK(CLK), .RN(RST_N), .Q(REG_B[11]), 
        .QN(N219) );
  DFFRX2TF \reg_B_reg[9]  ( .D(N454), .CK(CLK), .RN(RST_N), .Q(REG_B[9]), .QN(
        N217) );
  DFFRX2TF \reg_B_reg[8]  ( .D(N457), .CK(CLK), .RN(RST_N), .Q(REG_B[8]), .QN(
        N216) );
  DFFRX2TF \reg_A_reg[15]  ( .D(N5120), .CK(CLK), .RN(RST_N), .Q(REG_A[15]), 
        .QN(N267) );
  DFFRX2TF \reg_A_reg[13]  ( .D(N626), .CK(CLK), .RN(RST_N), .Q(REG_A[13]), 
        .QN(N277) );
  DFFRX2TF \reg_A_reg[11]  ( .D(N5130), .CK(CLK), .RN(RST_N), .Q(REG_A[11]), 
        .QN(N287) );
  DFFRX2TF \reg_A_reg[9]  ( .D(N610), .CK(CLK), .RN(RST_N), .Q(REG_A[9]), .QN(
        N266) );
  DFFRX2TF \reg_A_reg[8]  ( .D(N598), .CK(CLK), .RN(RST_N), .Q(REG_A[8]), .QN(
        N274) );
  DFFRX2TF \reg_A_reg[14]  ( .D(N634), .CK(CLK), .RN(RST_N), .Q(REG_A[14]), 
        .QN(N278) );
  DFFRX2TF \reg_A_reg[10]  ( .D(N5140), .CK(CLK), .RN(RST_N), .Q(REG_A[10]), 
        .QN(N283) );
  DFFRX2TF \reg_A_reg[12]  ( .D(N618), .CK(CLK), .RN(RST_N), .Q(REG_A[12]), 
        .QN(N276) );
  DFFRX2TF \reg_A_reg[6]  ( .D(N602), .CK(CLK), .RN(RST_N), .Q(REG_A[6]), .QN(
        N279) );
  DFFRX2TF \reg_A_reg[4]  ( .D(N606), .CK(CLK), .RN(RST_N), .Q(REG_A[4]), .QN(
        N280) );
  DFFNSRX2TF \id_ir_reg[4]  ( .D(N532), .CKN(CLK), .SN(1'b1), .RN(RST_N), .QN(
        N412) );
  DFFNSRX2TF \id_ir_reg[6]  ( .D(N536), .CKN(CLK), .SN(1'b1), .RN(RST_N), .QN(
        N411) );
  DFFNSRX2TF \gr_reg[1][7]  ( .D(N1074), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N794) );
  DFFNSRX2TF \gr_reg[1][6]  ( .D(N1075), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        IO_CONTROL[6]), .QN(N795) );
  DFFNSRX2TF \gr_reg[2][13]  ( .D(N1108), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N772) );
  DFFNSRX2TF \gr_reg[1][13]  ( .D(N1116), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N788) );
  DFFNSRX2TF \gr_reg[1][12]  ( .D(N1117), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N789) );
  DFFNSRX2TF \gr_reg[1][11]  ( .D(N1118), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N790) );
  DFFNSRX2TF \gr_reg[1][10]  ( .D(N1119), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N791) );
  DFFNSRX2TF \gr_reg[1][9]  ( .D(N1120), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N792) );
  DFFNSRX2TF \gr_reg[1][8]  ( .D(N1121), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N793) );
  DFFNSRX2TF \gr_reg[2][15]  ( .D(N1106), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N770) );
  DFFNSRX2TF \gr_reg[2][14]  ( .D(N1107), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N771) );
  DFFNSRX2TF \gr_reg[1][15]  ( .D(N1114), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N786) );
  DFFNSRX2TF \gr_reg[1][14]  ( .D(N1115), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N787) );
  DFFNSRX2TF \gr_reg[0][7]  ( .D(N1082), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N810) );
  DFFNSRX2TF \gr_reg[0][5]  ( .D(N1084), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N812) );
  DFFNSRX2TF \gr_reg[0][3]  ( .D(N1086), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N814) );
  DFFNSRX2TF \gr_reg[0][2]  ( .D(N1087), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N815) );
  DFFNSRX2TF \gr_reg[0][1]  ( .D(N1088), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N816) );
  DFFNSRX2TF \gr_reg[0][0]  ( .D(N1089), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N817) );
  DFFNSRX2TF \gr_reg[0][12]  ( .D(N1125), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N805) );
  DFFNSRX2TF \gr_reg[0][11]  ( .D(N1126), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N806) );
  DFFNSRX2TF \gr_reg[0][10]  ( .D(N1127), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N807) );
  DFFNSRX2TF \gr_reg[0][9]  ( .D(N1128), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N808) );
  DFFNSRX2TF \gr_reg[0][8]  ( .D(N1129), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N809) );
  DFFNSRX2TF \gr_reg[0][6]  ( .D(N1083), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N811) );
  DFFNSRX2TF \gr_reg[0][4]  ( .D(N1085), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N813) );
  DFFNSRX2TF \gr_reg[4][12]  ( .D(N1093), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N741) );
  DFFNSRX2TF \gr_reg[4][11]  ( .D(N1094), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N742) );
  DFFNSRX2TF \gr_reg[4][10]  ( .D(N1095), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N743) );
  DFFNSRX2TF \gr_reg[0][13]  ( .D(N1124), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N804) );
  DFFNSRX2TF \gr_reg[4][13]  ( .D(N1092), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N740) );
  DFFNSRX2TF \gr_reg[0][15]  ( .D(N1122), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N802) );
  DFFNSRX2TF \gr_reg[0][14]  ( .D(N1123), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N803) );
  DFFNSRX2TF \gr_reg[4][15]  ( .D(N1090), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N738) );
  DFFNSRX2TF \gr_reg[4][14]  ( .D(N1091), .CKN(CLK), .SN(1'b1), .RN(RST_N), 
        .QN(N739) );
  DFFNSRX2TF \id_ir_reg[11]  ( .D(N583), .CKN(CLK), .SN(1'b1), .RN(RST_N), .Q(
        N301), .QN(N53) );
  DFFSX2TF \reg_B_reg[1]  ( .D(N58), .CK(CLK), .SN(RST_N), .Q(N210), .QN(
        REG_B[1]) );
  NOR2X1TF U3 ( .A(N161), .B(N169), .Y(N580) );
  NAND3X1TF U4 ( .A(N169), .B(N426), .C(N934), .Y(N487) );
  AOI221X1TF U5 ( .A0(\SUB_X_276_4_B[0] ), .A1(N1014), .B0(N54), .B1(N59), 
        .C0(REG_B[1]), .Y(N694) );
  NAND2X1TF U6 ( .A(N961), .B(N954), .Y(N948) );
  NAND2X1TF U7 ( .A(N961), .B(N955), .Y(N950) );
  NOR2X1TF U8 ( .A(N896), .B(N917), .Y(N898) );
  NOR2X1TF U9 ( .A(N161), .B(CODE_TYPE[2]), .Y(N934) );
  NAND2X1TF U10 ( .A(CODE_TYPE[2]), .B(N580), .Y(N894) );
  NAND2X1TF U11 ( .A(N695), .B(N4670), .Y(N449) );
  NAND2X1TF U12 ( .A(N695), .B(N500), .Y(N497) );
  INVX2TF U13 ( .A(N1016), .Y(N1209) );
  OAI2BB1X1TF U14 ( .A0N(N202), .A1N(N514), .B0(N325), .Y(N1223) );
  NAND2X1TF U15 ( .A(STATE[1]), .B(IS_I_ADDR), .Y(N1142) );
  AOI211X1TF U16 ( .A0(N1640), .A1(N555), .B0(N554), .C0(N576), .Y(N574) );
  NAND2X1TF U17 ( .A(N936), .B(N937), .Y(N308) );
  NAND2X1TF U18 ( .A(STATE[1]), .B(STATE[2]), .Y(N523) );
  OAI2BB1X1TF U19 ( .A0N(N216), .A1N(N303), .B0(N674), .Y(N1) );
  AOI22X1TF U20 ( .A0(N420), .A1(N274), .B0(REG_A[8]), .B1(N295), .Y(N2) );
  AOI22X1TF U21 ( .A0(N670), .A1(N404), .B0(N159), .B1(N475), .Y(N3) );
  AOI32X1TF U22 ( .A0(N2), .A1(N3), .A2(N204), .B0(N216), .B1(N3), .Y(N4) );
  AOI222XLTF U23 ( .A0(N839), .A1(N851), .B0(N841), .B1(N1630), .C0(N671), 
        .C1(N406), .Y(N5) );
  AOI22X1TF U24 ( .A0(N669), .A1(N297), .B0(N509), .B1(N202), .Y(N6) );
  NAND2X1TF U25 ( .A(N5), .B(N6), .Y(N7) );
  AOI211X1TF U26 ( .A0(REG_A[8]), .A1(N1), .B0(N4), .C0(N7), .Y(N1178) );
  NAND2X1TF U27 ( .A(I_ADDR[2]), .B(I_ADDR[1]), .Y(N8) );
  AOI32X1TF U28 ( .A0(I_ADDR[2]), .A1(N572), .A2(I_ADDR[1]), .B0(N203), .B1(
        N572), .Y(N9) );
  AOI22XLTF U29 ( .A0(I_ADDR[3]), .A1(N9), .B0(D_ADDR[3]), .B1(N576), .Y(N10)
         );
  OAI31X1TF U30 ( .A0(N203), .A1(I_ADDR[3]), .A2(N8), .B0(N10), .Y(N657) );
  AOI22X1TF U31 ( .A0(REG_A[6]), .A1(N295), .B0(N303), .B1(N279), .Y(N11) );
  AOI21X1TF U32 ( .A0(N11), .A1(N204), .B0(N214), .Y(N12) );
  AOI222XLTF U33 ( .A0(N819), .A1(N1630), .B0(N875), .B1(N867), .C0(N406), 
        .C1(N870), .Y(N13) );
  OAI2BB1X1TF U34 ( .A0N(N214), .A1N(N303), .B0(N674), .Y(N14) );
  AOI222XLTF U35 ( .A0(N14), .A1(REG_A[6]), .B0(N473), .B1(N180), .C0(N650), 
        .C1(N851), .Y(N15) );
  NAND2X1TF U36 ( .A(N868), .B(N297), .Y(N16) );
  NAND3X1TF U37 ( .A(N13), .B(N15), .C(N16), .Y(N17) );
  AOI211X1TF U38 ( .A0(N202), .A1(N507), .B0(N12), .C0(N17), .Y(N1165) );
  AOI32X1TF U39 ( .A0(N563), .A1(N572), .A2(I_ADDR[4]), .B0(N578), .B1(N572), 
        .Y(N18) );
  AOI22XLTF U40 ( .A0(I_ADDR[5]), .A1(N18), .B0(D_ADDR[5]), .B1(N576), .Y(N19)
         );
  OAI31X1TF U41 ( .A0(N203), .A1(I_ADDR[5]), .A2(N562), .B0(N19), .Y(N659) );
  AOI22X1TF U42 ( .A0(REG_A[4]), .A1(N295), .B0(N303), .B1(N280), .Y(N20) );
  AOI21X1TF U43 ( .A0(N20), .A1(N204), .B0(N212), .Y(N21) );
  AOI222XLTF U44 ( .A0(N839), .A1(N714), .B0(N840), .B1(N1630), .C0(N670), 
        .C1(N406), .Y(N22) );
  OAI2BB1X1TF U45 ( .A0N(N212), .A1N(N303), .B0(N674), .Y(N23) );
  AOI222XLTF U46 ( .A0(N23), .A1(REG_A[4]), .B0(N159), .B1(N471), .C0(N841), 
        .C1(N851), .Y(N24) );
  NAND2X1TF U47 ( .A(N671), .B(N297), .Y(N25) );
  NAND3X1TF U48 ( .A(N22), .B(N24), .C(N25), .Y(N26) );
  AOI211X1TF U49 ( .A0(N874), .A1(N505), .B0(N21), .C0(N26), .Y(N1171) );
  CLKINVX1TF U50 ( .A(N559), .Y(N27) );
  OAI21X1TF U51 ( .A0(N578), .A1(I_ADDR[6]), .B0(N27), .Y(N28) );
  AOI22XLTF U52 ( .A0(I_ADDR[7]), .A1(N28), .B0(D_ADDR[7]), .B1(N576), .Y(N29)
         );
  OAI31X1TF U53 ( .A0(N203), .A1(I_ADDR[7]), .A2(N557), .B0(N29), .Y(N661) );
  AOI21X1TF U54 ( .A0(N302), .A1(N219), .B0(N876), .Y(N30) );
  OAI21X1TF U55 ( .A0(N879), .A1(REG_A[11]), .B0(N204), .Y(N31) );
  AOI21X1TF U56 ( .A0(REG_A[11]), .A1(N421), .B0(N31), .Y(N32) );
  CLKINVX1TF U57 ( .A(REG_B[11]), .Y(N33) );
  AOI22X1TF U58 ( .A0(N297), .A1(N706), .B0(N406), .B1(N860), .Y(N34) );
  CLKINVX1TF U59 ( .A(N857), .Y(N35) );
  AOI222XLTF U60 ( .A0(N35), .A1(N851), .B0(N850), .B1(N1630), .C0(N854), .C1(
        N404), .Y(N36) );
  OAI211X1TF U61 ( .A0(N32), .A1(N33), .B0(N34), .C0(N36), .Y(N37) );
  AOI21X1TF U62 ( .A0(N202), .A1(N512), .B0(N37), .Y(N38) );
  NAND2X1TF U63 ( .A(N159), .B(N478), .Y(N39) );
  OAI211X1TF U64 ( .A0(N287), .A1(N30), .B0(N38), .C0(N39), .Y(N1196) );
  NOR2X1TF U65 ( .A(N752), .B(N196), .Y(N40) );
  OAI22X1TF U66 ( .A0(N784), .A1(N193), .B0(N816), .B1(N170), .Y(N41) );
  OAI22X1TF U67 ( .A0(N1218), .A1(N261), .B0(N768), .B1(N1227), .Y(N42) );
  OAI22X1TF U68 ( .A0(N210), .A1(N1236), .B0(N800), .B1(N182), .Y(N43) );
  NOR4XLTF U69 ( .A(N40), .B(N41), .C(N42), .D(N43), .Y(N58) );
  AOI22XLTF U70 ( .A0(N576), .A1(D_ADDR[1]), .B0(I_ADDR[1]), .B1(N574), .Y(N44) );
  OAI21X1TF U71 ( .A0(I_ADDR[1]), .A1(N203), .B0(N44), .Y(N654) );
  AOI21X1TF U72 ( .A0(N56), .A1(REG_A[9]), .B0(N646), .Y(N45) );
  NAND3X1TF U73 ( .A(N612), .B(N615), .C(N45), .Y(N819) );
  NOR2BX1TF U74 ( .AN(N424), .B(N938), .Y(N416) );
  OAI22X1TF U75 ( .A0(N775), .A1(N193), .B0(N807), .B1(N170), .Y(N46) );
  OAI22X1TF U76 ( .A0(N791), .A1(N181), .B0(N743), .B1(N195), .Y(N47) );
  OAI22X1TF U77 ( .A0(N1226), .A1(N269), .B0(N201), .B1(N759), .Y(N48) );
  NOR3X1TF U78 ( .A(N46), .B(N47), .C(N48), .Y(N49) );
  OAI21X1TF U79 ( .A0(N218), .A1(N1236), .B0(N49), .Y(N5110) );
  OAI22X1TF U80 ( .A0(N160), .A1(N1014), .B0(N801), .B1(N173), .Y(N50) );
  AOI22X1TF U81 ( .A0(IO_OFFSET[0]), .A1(N1016), .B0(N1015), .B1(
        IO_DATAOUTA[0]), .Y(N51) );
  OAI21X1TF U82 ( .A0(N177), .A1(N817), .B0(N51), .Y(N52) );
  AOI211X1TF U83 ( .A0(N175), .A1(IO_DATAOUTB[0]), .B0(N50), .C0(N52), .Y(N97)
         );
  MX2X4TF U84 ( .A(ADD_X_276_3_N18), .B(ADD_X_276_3_N17), .S0(ADD_X_276_3_N21), 
        .Y(ADD_X_276_3_N16) );
  ADDFHX2TF U85 ( .A(N210), .B(REG_A[1]), .CI(SUB_X_276_4_N16), .CO(
        SUB_X_276_4_N15), .S(N502) );
  NAND2BX2TF U86 ( .AN(REG_A[0]), .B(\SUB_X_276_4_B[0] ), .Y(SUB_X_276_4_N16)
         );
  BUFX4TF U87 ( .A(REG_B[0]), .Y(\SUB_X_276_4_B[0] ) );
  AND2X2TF U88 ( .A(REG_B[1]), .B(\SUB_X_276_4_B[0] ), .Y(N56) );
  INVX2TF U89 ( .A(N289), .Y(N161) );
  NAND2X1TF U90 ( .A(IS_I_ADDR), .B(N270), .Y(N1137) );
  INVXLTF U91 ( .A(REG_B[3]), .Y(N60) );
  AOI22XLTF U92 ( .A0(N444), .A1(N4760), .B0(N787), .B1(N443), .Y(N1115) );
  OAI22XLTF U93 ( .A0(N739), .A1(N195), .B0(N787), .B1(N181), .Y(N901) );
  AOI22XLTF U94 ( .A0(N444), .A1(N4820), .B0(N786), .B1(N443), .Y(N1114) );
  OAI22XLTF U95 ( .A0(N738), .A1(N195), .B0(N786), .B1(N181), .Y(N1232) );
  OAI22XLTF U96 ( .A0(N803), .A1(N209), .B0(N771), .B1(N192), .Y(N1029) );
  OAI22XLTF U97 ( .A0(N771), .A1(N1210), .B0(N1209), .B1(N739), .Y(N1211) );
  OAI22XLTF U98 ( .A0(N803), .A1(N171), .B0(N771), .B1(N194), .Y(N902) );
  OAI22XLTF U99 ( .A0(N802), .A1(N208), .B0(N770), .B1(N191), .Y(N1026) );
  OAI22XLTF U100 ( .A0(N770), .A1(N1210), .B0(N1209), .B1(N738), .Y(N1017) );
  OAI22XLTF U101 ( .A0(N802), .A1(N171), .B0(N770), .B1(N194), .Y(N1233) );
  AOI22XLTF U102 ( .A0(N444), .A1(N4700), .B0(N791), .B1(N443), .Y(N1119) );
  AOI22XLTF U103 ( .A0(N444), .A1(N4710), .B0(N790), .B1(N443), .Y(N1118) );
  OAI22XLTF U104 ( .A0(N742), .A1(N195), .B0(N790), .B1(N181), .Y(N1192) );
  AOI22XLTF U105 ( .A0(N444), .A1(N4720), .B0(N789), .B1(N443), .Y(N1117) );
  OAI22XLTF U106 ( .A0(N741), .A1(N195), .B0(N789), .B1(N181), .Y(N909) );
  AOI22XLTF U107 ( .A0(N444), .A1(N4740), .B0(N788), .B1(N443), .Y(N1116) );
  OAI22XLTF U108 ( .A0(N740), .A1(N195), .B0(N788), .B1(N181), .Y(N905) );
  OAI22XLTF U109 ( .A0(N804), .A1(N208), .B0(N772), .B1(N191), .Y(N1032) );
  OAI22XLTF U110 ( .A0(N772), .A1(N1210), .B0(N1209), .B1(N740), .Y(N1199) );
  OAI22XLTF U111 ( .A0(N804), .A1(N171), .B0(N772), .B1(N193), .Y(N906) );
  AOI22XLTF U112 ( .A0(N494), .A1(N5070), .B0(N795), .B1(N493), .Y(N1075) );
  AOI22XLTF U113 ( .A0(N494), .A1(N5090), .B0(N794), .B1(N493), .Y(N1074) );
  AOI31XLTF U114 ( .A0(N411), .A1(N412), .A2(N945), .B0(N944), .Y(N1215) );
  AO21X4TF U115 ( .A0(N482), .A1(N159), .B0(N356), .Y(N357) );
  AOI211X1TF U167 ( .A0(REG_B[1]), .A1(N700), .B0(N699), .C0(N698), .Y(N702)
         );
  INVX2TF U168 ( .A(N179), .Y(N159) );
  OA22X1TF U169 ( .A0(N412), .A1(N949), .B0(N962), .B1(N948), .Y(N1213) );
  INVX1TF U170 ( .A(N409), .Y(N887) );
  CLKINVX2TF U171 ( .A(N404), .Y(N662) );
  INVX2TF U172 ( .A(N956), .Y(N160) );
  AND4X1TF U173 ( .A(N261), .B(N259), .C(N269), .D(N898), .Y(N1229) );
  NAND2BXLTF U174 ( .AN(N960), .B(N423), .Y(N307) );
  OAI21XLTF U175 ( .A0(N893), .A1(N161), .B0(N311), .Y(N312) );
  CLKINVX1TF U176 ( .A(N558), .Y(N561) );
  NAND3XLTF U177 ( .A(N161), .B(N940), .C(N426), .Y(N431) );
  NAND2X1TF U178 ( .A(N161), .B(N55), .Y(N938) );
  NAND2XLTF U179 ( .A(D_WE), .B(N544), .Y(N436) );
  OAI22X1TF U180 ( .A0(N813), .A1(N208), .B0(N781), .B1(N191), .Y(N988) );
  OAI22X1TF U181 ( .A0(N807), .A1(N208), .B0(N775), .B1(N191), .Y(N1041) );
  OAI22X1TF U182 ( .A0(N810), .A1(N208), .B0(N778), .B1(N191), .Y(N966) );
  OAI22X1TF U183 ( .A0(N817), .A1(N208), .B0(N785), .B1(N191), .Y(N1011) );
  OAI22X1TF U184 ( .A0(N815), .A1(N170), .B0(N783), .B1(N193), .Y(N1147) );
  OAI22X1TF U185 ( .A0(N744), .A1(N195), .B0(N792), .B1(N181), .Y(N913) );
  OAI22X1TF U186 ( .A0(N745), .A1(N195), .B0(N793), .B1(N181), .Y(N926) );
  OAI22X1TF U187 ( .A0(N812), .A1(N170), .B0(N780), .B1(N193), .Y(N976) );
  OAI22X1TF U188 ( .A0(N814), .A1(N170), .B0(N782), .B1(N193), .Y(N1180) );
  OAI22X1TF U189 ( .A0(N813), .A1(N170), .B0(N781), .B1(N193), .Y(N919) );
  AOI22X1TF U190 ( .A0(N494), .A1(N5040), .B0(N798), .B1(N493), .Y(N1078) );
  AOI22X1TF U191 ( .A0(N496), .A1(N5050), .B0(N781), .B1(N495), .Y(N1069) );
  AOI22X1TF U192 ( .A0(N444), .A1(N4690), .B0(N792), .B1(N443), .Y(N1120) );
  AOI22X1TF U193 ( .A0(N447), .A1(N4710), .B0(N774), .B1(N445), .Y(N1110) );
  AOI22X1TF U194 ( .A0(N494), .A1(N5060), .B0(N796), .B1(N493), .Y(N1076) );
  AOI22X1TF U195 ( .A0(N494), .A1(N5020), .B0(N800), .B1(N493), .Y(N1080) );
  AOI22X1TF U196 ( .A0(N499), .A1(N5090), .B0(N762), .B1(N498), .Y(N1058) );
  AOI22X1TF U197 ( .A0(N496), .A1(N5040), .B0(N782), .B1(N495), .Y(N1070) );
  AOI22X1TF U198 ( .A0(N447), .A1(N4720), .B0(N773), .B1(N445), .Y(N1109) );
  AOI22X1TF U199 ( .A0(N447), .A1(N4700), .B0(N775), .B1(N445), .Y(N1111) );
  AOI22X1TF U200 ( .A0(N447), .A1(N4690), .B0(N776), .B1(N445), .Y(N1112) );
  AOI22X1TF U201 ( .A0(N499), .A1(N5070), .B0(N763), .B1(N498), .Y(N1059) );
  AOI22X1TF U202 ( .A0(N462), .A1(N4680), .B0(N761), .B1(N461), .Y(N1105) );
  AOI22X1TF U203 ( .A0(N462), .A1(N4700), .B0(N759), .B1(N461), .Y(N1103) );
  AOI22X1TF U204 ( .A0(N499), .A1(N5010), .B0(N769), .B1(N498), .Y(N1065) );
  AOI22X1TF U205 ( .A0(N499), .A1(N5020), .B0(N768), .B1(N498), .Y(N1064) );
  AOI22X1TF U206 ( .A0(N462), .A1(N4710), .B0(N758), .B1(N461), .Y(N1102) );
  AOI22X1TF U207 ( .A0(N496), .A1(N5010), .B0(N785), .B1(N495), .Y(N1073) );
  AOI22X1TF U208 ( .A0(N447), .A1(N4680), .B0(N777), .B1(N445), .Y(N1113) );
  AOI22X1TF U209 ( .A0(N499), .A1(N5030), .B0(N767), .B1(N498), .Y(N1063) );
  AOI22X1TF U210 ( .A0(N496), .A1(N5090), .B0(N778), .B1(N495), .Y(N1066) );
  AOI22X1TF U211 ( .A0(N462), .A1(N4720), .B0(N757), .B1(N461), .Y(N1101) );
  AOI22X1TF U212 ( .A0(N496), .A1(N5070), .B0(N779), .B1(N495), .Y(N1067) );
  AOI22X1TF U213 ( .A0(N462), .A1(N4690), .B0(N760), .B1(N461), .Y(N1104) );
  AND2X2TF U214 ( .A(N964), .B(N187), .Y(N207) );
  AND2X2TF U215 ( .A(N965), .B(N187), .Y(N1049) );
  AND2X2TF U216 ( .A(N187), .B(N265), .Y(N1136) );
  NAND2XLTF U217 ( .A(N591), .B(N433), .Y(N585) );
  INVX2TF U218 ( .A(N827), .Y(N162) );
  AND2X2TF U219 ( .A(OPER3_R3[0]), .B(N900), .Y(N1230) );
  AO22X1TF U220 ( .A0(N963), .A1(N952), .B0(N413), .B1(N951), .Y(N1208) );
  OAI211X1TF U221 ( .A0(STATE[1]), .A1(N533), .B0(N531), .C0(N544), .Y(
        NEXT_STATE[0]) );
  INVX2TF U222 ( .A(N186), .Y(N187) );
  AND2X2TF U223 ( .A(OPER3_R3[1]), .B(N897), .Y(N1228) );
  OA21X2TF U224 ( .A0(N891), .A1(N308), .B0(N410), .Y(N409) );
  OAI2BB1X1TF U225 ( .A0N(N314), .A1N(N941), .B0(N313), .Y(N371) );
  AND2X2TF U226 ( .A(N898), .B(OPER3_R3[2]), .Y(N1231) );
  NAND3X2TF U227 ( .A(N898), .B(OPER3_R3[0]), .C(OPER3_R3[1]), .Y(N1227) );
  NAND2XLTF U228 ( .A(N184), .B(REG_A[3]), .Y(N691) );
  CLKAND2X2TF U229 ( .A(N426), .B(N550), .Y(N408) );
  CLKAND2X2TF U230 ( .A(N383), .B(N550), .Y(N394) );
  INVX1TF U231 ( .A(N422), .Y(N382) );
  INVX1TF U232 ( .A(N582), .Y(N310) );
  OR2X1TF U233 ( .A(CODE_TYPE[3]), .B(N582), .Y(N971) );
  INVX2TF U234 ( .A(N1137), .Y(N189) );
  INVX2TF U235 ( .A(N56), .Y(N1650) );
  NOR2X1TF U236 ( .A(N260), .B(N696), .Y(N965) );
  INVX2TF U237 ( .A(N827), .Y(N1630) );
  CLKBUFX2TF U238 ( .A(N556), .Y(N1640) );
  NOR3X1TF U239 ( .A(N679), .B(N262), .C(N523), .Y(N556) );
  INVX2TF U240 ( .A(N56), .Y(N166) );
  INVX2TF U241 ( .A(N1142), .Y(N167) );
  INVX2TF U242 ( .A(N1142), .Y(N168) );
  INVX2TF U243 ( .A(N301), .Y(N169) );
  INVX2TF U244 ( .A(N1229), .Y(N170) );
  INVX2TF U245 ( .A(N1229), .Y(N171) );
  INVX2TF U246 ( .A(N1208), .Y(N172) );
  INVX2TF U247 ( .A(N1208), .Y(N173) );
  INVX2TF U248 ( .A(N1213), .Y(N174) );
  INVX2TF U249 ( .A(N1213), .Y(N175) );
  INVX2TF U250 ( .A(N1215), .Y(N176) );
  INVX2TF U251 ( .A(N176), .Y(N177) );
  INVX2TF U252 ( .A(N176), .Y(N178) );
  INVX2TF U253 ( .A(N371), .Y(N179) );
  INVX2TF U254 ( .A(N179), .Y(N180) );
  INVX2TF U255 ( .A(N1230), .Y(N181) );
  INVX2TF U256 ( .A(N1230), .Y(N182) );
  INVX2TF U257 ( .A(N843), .Y(N183) );
  INVX2TF U258 ( .A(N843), .Y(N184) );
  INVX2TF U259 ( .A(N1048), .Y(N186) );
  INVX2TF U260 ( .A(N186), .Y(N188) );
  NOR3X2TF U261 ( .A(N260), .B(N275), .C(N265), .Y(N964) );
  AOI22X2TF U262 ( .A0(N1640), .A1(D_ADDR[8]), .B0(D_DATAIN[7]), .B1(N543), 
        .Y(N5090) );
  AOI22X2TF U263 ( .A0(N1640), .A1(D_ADDR[7]), .B0(D_DATAIN[6]), .B1(N543), 
        .Y(N5070) );
  AOI22X2TF U264 ( .A0(D_ADDR[1]), .A1(N1640), .B0(D_DATAIN[0]), .B1(N543), 
        .Y(N5010) );
  AOI22X2TF U265 ( .A0(N1640), .A1(D_ADDR[5]), .B0(D_DATAIN[4]), .B1(N543), 
        .Y(N5050) );
  AOI22X2TF U266 ( .A0(N1640), .A1(D_ADDR[3]), .B0(D_DATAIN[2]), .B1(N543), 
        .Y(N5030) );
  AOI22X2TF U267 ( .A0(N1640), .A1(D_ADDR[2]), .B0(D_DATAIN[1]), .B1(N543), 
        .Y(N5020) );
  AOI22X2TF U268 ( .A0(N1640), .A1(D_ADDR[4]), .B0(D_DATAIN[3]), .B1(N543), 
        .Y(N5040) );
  AOI2BB2X2TF U269 ( .B0(D_DATAIN[4]), .B1(N439), .A0N(N418), .A1N(N488), .Y(
        N4720) );
  AOI2BB2X2TF U270 ( .B0(D_DATAIN[0]), .B1(N439), .A0N(N425), .A1N(N488), .Y(
        N4680) );
  AOI2BB2X2TF U271 ( .B0(D_DATAIN[3]), .B1(N439), .A0N(N415), .A1N(N488), .Y(
        N4710) );
  AOI2BB2X2TF U272 ( .B0(D_DATAIN[2]), .B1(N439), .A0N(N427), .A1N(N488), .Y(
        N4700) );
  AOI22X2TF U273 ( .A0(N1640), .A1(D_ADDR[6]), .B0(D_DATAIN[5]), .B1(N543), 
        .Y(N5060) );
  AOI22X2TF U274 ( .A0(REG_C[15]), .A1(N440), .B0(N439), .B1(D_DATAIN[7]), .Y(
        N4820) );
  AOI22X2TF U275 ( .A0(REG_C[14]), .A1(N440), .B0(N439), .B1(D_DATAIN[6]), .Y(
        N4760) );
  AOI2BB2X2TF U276 ( .B0(D_DATAIN[5]), .B1(N439), .A0N(N414), .A1N(N488), .Y(
        N4740) );
  NOR3X4TF U277 ( .A(N697), .B(N696), .C(N449), .Y(N462) );
  NOR3X4TF U278 ( .A(N697), .B(N696), .C(N497), .Y(N499) );
  NOR3X4TF U279 ( .A(N696), .B(N260), .C(N497), .Y(N496) );
  INVX2TF U280 ( .A(N1137), .Y(N190) );
  INVX2TF U281 ( .A(N1049), .Y(N191) );
  INVX2TF U282 ( .A(N1049), .Y(N192) );
  INVX2TF U283 ( .A(N1228), .Y(N193) );
  INVX2TF U284 ( .A(N1228), .Y(N194) );
  INVX2TF U285 ( .A(N1231), .Y(N195) );
  INVX2TF U286 ( .A(N1231), .Y(N196) );
  INVX2TF U287 ( .A(N1136), .Y(N197) );
  INVX2TF U288 ( .A(N1136), .Y(N198) );
  CLKBUFX2TF U289 ( .A(N398), .Y(N199) );
  CLKBUFX2TF U290 ( .A(N1134), .Y(N200) );
  NOR2BX2TF U291 ( .AN(N188), .B(N962), .Y(N1134) );
  CLKBUFX2TF U292 ( .A(N1227), .Y(N201) );
  CLKBUFX2TF U293 ( .A(N160), .Y(N300) );
  NAND2X1TF U294 ( .A(N210), .B(N54), .Y(N675) );
  INVX2TF U295 ( .A(N675), .Y(N862) );
  CLKBUFX2TF U296 ( .A(N874), .Y(N202) );
  AOI21X2TF U297 ( .A0(N513), .A1(N202), .B0(N363), .Y(N400) );
  NAND2X2TF U298 ( .A(N307), .B(N306), .Y(N874) );
  OAI221X1TF U299 ( .A0(\SUB_X_276_4_B[0] ), .A1(REG_A[14]), .B0(N54), .B1(
        REG_A[15]), .C0(N210), .Y(N652) );
  OAI21XLTF U300 ( .A0(N675), .A1(N821), .B0(N674), .Y(N683) );
  OAI21XLTF U301 ( .A0(N970), .A1(N894), .B0(N674), .Y(N432) );
  NOR2X2TF U302 ( .A(N57), .B(N211), .Y(N869) );
  NOR3X2TF U303 ( .A(STATE[2]), .B(STATE[3]), .C(N679), .Y(IS_I_ADDR) );
  AOI2BB2X2TF U304 ( .B0(D_DATAIN[1]), .B1(N439), .A0N(N419), .A1N(N488), .Y(
        N4690) );
  INVX2TF U305 ( .A(N569), .Y(N203) );
  NAND2X1TF U306 ( .A(N556), .B(N552), .Y(N578) );
  NOR3X4TF U307 ( .A(N296), .B(N969), .C(N382), .Y(N395) );
  INVX2TF U308 ( .A(N881), .Y(N204) );
  NOR2BX1TF U309 ( .AN(N591), .B(N953), .Y(N838) );
  CLKBUFX2TF U310 ( .A(N1047), .Y(N205) );
  CLKBUFX2TF U311 ( .A(N1236), .Y(N206) );
  OAI21X2TF U312 ( .A0(N895), .A1(N917), .B0(N961), .Y(N1218) );
  INVX2TF U313 ( .A(N207), .Y(N208) );
  INVX2TF U314 ( .A(N207), .Y(N209) );
  NOR3X4TF U315 ( .A(N696), .B(N260), .C(N449), .Y(N447) );
  XOR2X1TF U316 ( .A(REG_A[0]), .B(\SUB_X_276_4_B[0] ), .Y(N501) );
  INVX2TF U317 ( .A(SUB_X_276_4_N1), .Y(N517) );
  ADDFHX2TF U318 ( .A(N223), .B(REG_A[15]), .CI(SUB_X_276_4_N2), .CO(
        SUB_X_276_4_N1), .S(N516) );
  OAI21X2TF U319 ( .A0(N390), .A1(N1224), .B0(N389), .Y(N641) );
  XOR2X2TF U320 ( .A(N393), .B(N385), .Y(N390) );
  XOR2X4TF U321 ( .A(N1223), .B(N384), .Y(N385) );
  OAI211XLTF U322 ( .A0(N393), .A1(N1225), .B0(N392), .C0(N391), .Y(N645) );
  AOI21X1TF U323 ( .A0(N487), .A1(N488), .B0(N553), .Y(N4670) );
  NAND3X2TF U324 ( .A(N896), .B(N1226), .C(N1218), .Y(N1236) );
  CLKXOR2X2TF U325 ( .A(N400), .B(N401), .Y(N384) );
  NAND2X2TF U326 ( .A(N963), .B(N187), .Y(N1047) );
  OAI22X1TF U327 ( .A0(N553), .A1(N488), .B0(N487), .B1(N489), .Y(N500) );
  AOI32XLTF U328 ( .A0(N169), .A1(N693), .A2(NF), .B0(N546), .B1(N161), .Y(
        N547) );
  NAND2X1TF U329 ( .A(CODE_TYPE[2]), .B(N169), .Y(N590) );
  NOR2X2TF U330 ( .A(STATE[3]), .B(N890), .Y(N961) );
  CLKBUFX2TF U331 ( .A(N1238), .Y(N296) );
  CLKBUFX2TF U332 ( .A(N676), .Y(N299) );
  NAND2X1TF U333 ( .A(N424), .B(N550), .Y(N674) );
  NOR2X1TF U334 ( .A(N161), .B(N590), .Y(N550) );
  NAND2X1TF U335 ( .A(N434), .B(N262), .Y(N489) );
  INVX2TF U336 ( .A(N556), .Y(N553) );
  AO21X1TF U337 ( .A0(N396), .A1(N1207), .B0(N1206), .Y(N633) );
  INVX2TF U338 ( .A(N948), .Y(N952) );
  OAI211X1TF U339 ( .A0(N943), .A1(N970), .B0(N942), .C0(N941), .Y(N954) );
  NAND2BX1TF U340 ( .AN(N938), .B(N53), .Y(N943) );
  NOR2X2TF U341 ( .A(CODE_TYPE[3]), .B(CODE_TYPE[4]), .Y(N426) );
  NAND2X1TF U342 ( .A(CODE_TYPE[3]), .B(CODE_TYPE[4]), .Y(N893) );
  OAI32X1TF U343 ( .A0(N1238), .A1(N960), .A2(N969), .B0(N410), .B1(N436), .Y(
        N1130) );
  NOR3BX1TF U344 ( .AN(N961), .B(N960), .C(N969), .Y(N1048) );
  NOR2X2TF U345 ( .A(N492), .B(N497), .Y(N494) );
  OAI211X1TF U346 ( .A0(N940), .A1(N937), .B0(N936), .C0(N935), .Y(N955) );
  NOR4X1TF U347 ( .A(N1237), .B(N1223), .C(N1196), .D(N378), .Y(N379) );
  AOI222XLTF U348 ( .A0(N832), .A1(N867), .B0(N689), .B1(N428), .C0(N831), 
        .C1(N869), .Y(N703) );
  OAI2BB1X2TF U349 ( .A0N(N202), .A1N(N515), .B0(N321), .Y(N1237) );
  OAI211X1TF U350 ( .A0(N263), .A1(N894), .B0(N893), .C0(N892), .Y(N917) );
  NAND3X1TF U351 ( .A(STATE[1]), .B(N679), .C(N268), .Y(N890) );
  NAND2X1TF U352 ( .A(N679), .B(N262), .Y(N551) );
  INVX2TF U353 ( .A(N590), .Y(N429) );
  NOR2X2TF U354 ( .A(CODE_TYPE[2]), .B(N169), .Y(N940) );
  NOR2X2TF U355 ( .A(N492), .B(N449), .Y(N444) );
  INVX2TF U356 ( .A(N4790), .Y(N485) );
  INVX2TF U357 ( .A(N487), .Y(N439) );
  INVX2TF U358 ( .A(N5080), .Y(N5100) );
  INVX2TF U359 ( .A(N489), .Y(N543) );
  NOR2X1TF U360 ( .A(N679), .B(N523), .Y(N434) );
  CLKBUFX2TF U361 ( .A(N397), .Y(N298) );
  NOR2X1TF U362 ( .A(N275), .B(N697), .Y(N963) );
  NOR2X2TF U363 ( .A(N296), .B(N381), .Y(N396) );
  AOI222X1TF U364 ( .A0(N841), .A1(N867), .B0(N840), .B1(N428), .C0(N839), 
        .C1(N869), .Y(N849) );
  NOR2X1TF U365 ( .A(N296), .B(N970), .Y(N383) );
  INVX2TF U366 ( .A(N395), .Y(N1224) );
  OR2X2TF U367 ( .A(N551), .B(N523), .Y(N1238) );
  INVX2TF U368 ( .A(N441), .Y(N442) );
  INVX2TF U369 ( .A(N490), .Y(N491) );
  NOR4BX1TF U370 ( .AN(START), .B(STATE[1]), .C(STATE[2]), .D(N551), .Y(N554)
         );
  INVX2TF U371 ( .A(N396), .Y(N1225) );
  AND2X2TF U372 ( .A(N383), .B(N380), .Y(N397) );
  AOI21X4TF U373 ( .A0(N516), .A1(N202), .B0(N357), .Y(N393) );
  AND2X2TF U374 ( .A(N264), .B(CODE_TYPE[4]), .Y(N423) );
  OR2X2TF U375 ( .A(N161), .B(N305), .Y(N960) );
  NOR4XLTF U376 ( .A(N421), .B(N303), .C(N416), .D(N202), .Y(N433) );
  OAI2BB1X1TF U377 ( .A0N(N523), .A1N(STATE[3]), .B0(N430), .Y(N163) );
  AOI31XLTF U378 ( .A0(N679), .A1(START), .A2(N545), .B0(N1640), .Y(N430) );
  AO22X1TF U379 ( .A0(N483), .A1(N416), .B0(N517), .B1(N202), .Y(N586) );
  OR3X1TF U380 ( .A(N190), .B(N435), .C(N529), .Y(N1131) );
  AOI211XLTF U381 ( .A0(N262), .A1(N890), .B0(N434), .C0(N288), .Y(N435) );
  AO22X1TF U382 ( .A0(N409), .A1(CF_BUF), .B0(N887), .B1(CF), .Y(N446) );
  AOI31XLTF U383 ( .A0(N693), .A1(N940), .A2(N426), .B0(N553), .Y(N525) );
  OAI2BB2XLTF U384 ( .B0(N189), .B1(N261), .A0N(N189), .A1N(I_DATAIN[1]), .Y(
        N526) );
  OAI2BB2XLTF U385 ( .B0(N189), .B1(N269), .A0N(N190), .A1N(I_DATAIN[2]), .Y(
        N528) );
  OAI2BB2XLTF U386 ( .B0(N190), .B1(N259), .A0N(N190), .A1N(I_DATAIN[0]), .Y(
        N524) );
  OAI2BB2XLTF U387 ( .B0(N189), .B1(N413), .A0N(N190), .A1N(I_DATAIN[5]), .Y(
        N534) );
  OAI2BB2XLTF U388 ( .B0(N190), .B1(N412), .A0N(N190), .A1N(I_DATAIN[4]), .Y(
        N532) );
  OAI2BB2XLTF U389 ( .B0(N167), .B1(N696), .A0N(N167), .A1N(I_DATAIN[1]), .Y(
        N587) );
  OAI2BB2XLTF U390 ( .B0(N168), .B1(N55), .A0N(N168), .A1N(I_DATAIN[5]), .Y(
        N579) );
  OAI2BB2XLTF U391 ( .B0(N167), .B1(N697), .A0N(N167), .A1N(I_DATAIN[0]), .Y(
        N589) );
  OAI2BB2XLTF U392 ( .B0(N167), .B1(N695), .A0N(N167), .A1N(I_DATAIN[2]), .Y(
        N5850) );
  OAI2BB2XLTF U393 ( .B0(N168), .B1(N693), .A0N(N168), .A1N(I_DATAIN[4]), .Y(
        N581) );
  INVX2TF U394 ( .A(N444), .Y(N443) );
  INVX2TF U395 ( .A(N462), .Y(N461) );
  INVX2TF U396 ( .A(N447), .Y(N445) );
  INVX2TF U397 ( .A(N496), .Y(N495) );
  INVX2TF U398 ( .A(N499), .Y(N498) );
  NAND2X1TF U399 ( .A(N570), .B(I_ADDR[8]), .Y(N555) );
  NOR3X1TF U400 ( .A(N376), .B(N1207), .C(N1156), .Y(N377) );
  INVX2TF U401 ( .A(N296), .Y(N410) );
  NAND2X1TF U402 ( .A(N347), .B(REG_A[15]), .Y(N857) );
  NAND2X2TF U403 ( .A(N210), .B(\SUB_X_276_4_B[0] ), .Y(N842) );
  NAND2X2TF U404 ( .A(N54), .B(REG_B[1]), .Y(N843) );
  NOR2X1TF U405 ( .A(N553), .B(N431), .Y(N164) );
  OAI21X1TF U406 ( .A0(N545), .A1(N537), .B0(N535), .Y(NEXT_STATE[1]) );
  OAI21X1TF U407 ( .A0(N268), .A1(N291), .B0(N262), .Y(N537) );
  AOI22X1TF U408 ( .A0(I_ADDR[0]), .A1(N720), .B0(N728), .B1(N288), .Y(
        D_DATAOUT[7]) );
  AOI22X1TF U409 ( .A0(I_ADDR[0]), .A1(N721), .B0(N729), .B1(N288), .Y(
        D_DATAOUT[6]) );
  AOI22X1TF U410 ( .A0(I_ADDR[0]), .A1(N722), .B0(N730), .B1(N288), .Y(
        D_DATAOUT[5]) );
  AOI22X1TF U411 ( .A0(I_ADDR[0]), .A1(N723), .B0(N731), .B1(N288), .Y(
        D_DATAOUT[4]) );
  AOI22X1TF U412 ( .A0(I_ADDR[0]), .A1(N724), .B0(N732), .B1(N288), .Y(
        D_DATAOUT[3]) );
  AOI22X1TF U413 ( .A0(I_ADDR[0]), .A1(N725), .B0(N733), .B1(N288), .Y(
        D_DATAOUT[2]) );
  AOI22X1TF U414 ( .A0(I_ADDR[0]), .A1(N726), .B0(N734), .B1(N288), .Y(
        D_DATAOUT[1]) );
  AOI22X1TF U415 ( .A0(I_ADDR[0]), .A1(N727), .B0(N735), .B1(N288), .Y(
        D_DATAOUT[0]) );
  OAI211X1TF U416 ( .A0(N545), .A1(N551), .B0(N651), .C0(N544), .Y(
        NEXT_STATE[2]) );
  OAI32X1TF U417 ( .A0(N543), .A1(N542), .A2(N541), .B0(N540), .B1(N543), .Y(
        N651) );
  NOR2X1TF U418 ( .A(N539), .B(N1137), .Y(N541) );
  NOR2X1TF U419 ( .A(STATE[1]), .B(STATE[2]), .Y(N545) );
  AOI211X1TF U420 ( .A0(N190), .A1(N539), .B0(N529), .C0(N527), .Y(N531) );
  NOR2X1TF U421 ( .A(N189), .B(N542), .Y(N535) );
  NOR3X1TF U422 ( .A(N523), .B(N262), .C(N291), .Y(N542) );
  NOR2X1TF U423 ( .A(IO_STATUS[0]), .B(IO_STATUS[1]), .Y(N540) );
  OAI31X1TF U424 ( .A0(STATE[1]), .A1(N268), .A2(N551), .B0(N489), .Y(N529) );
  OAI21X1TF U425 ( .A0(N753), .A1(N197), .B0(N1013), .Y(N486) );
  AOI211X1TF U426 ( .A0(N1134), .A1(IO_DATAOUTB[0]), .B0(N1012), .C0(N1011), 
        .Y(N1013) );
  OAI22X1TF U427 ( .A0(N188), .A1(N735), .B0(N801), .B1(N1047), .Y(N1012) );
  OAI21X1TF U428 ( .A0(N743), .A1(N197), .B0(N1043), .Y(N520) );
  AOI211X1TF U429 ( .A0(N1134), .A1(IO_DATAOUTB[10]), .B0(N1042), .C0(N1041), 
        .Y(N1043) );
  OAI22X1TF U430 ( .A0(N187), .A1(N725), .B0(N791), .B1(N1047), .Y(N1042) );
  OAI21X1TF U431 ( .A0(N740), .A1(N197), .B0(N1034), .Y(N5170) );
  AOI211X1TF U432 ( .A0(N1134), .A1(N285), .B0(N1033), .C0(N1032), .Y(N1034)
         );
  OAI22X1TF U433 ( .A0(N188), .A1(N722), .B0(N788), .B1(N1047), .Y(N1033) );
  OAI21X1TF U434 ( .A0(N749), .A1(N197), .B0(N990), .Y(N4750) );
  AOI211X1TF U435 ( .A0(N1134), .A1(IO_DATAOUTB[4]), .B0(N989), .C0(N988), .Y(
        N990) );
  OAI22X1TF U436 ( .A0(N187), .A1(N731), .B0(N797), .B1(N1047), .Y(N989) );
  OAI21X1TF U437 ( .A0(N746), .A1(N197), .B0(N968), .Y(N460) );
  AOI211X1TF U438 ( .A0(N1134), .A1(IO_DATAOUTB[7]), .B0(N967), .C0(N966), .Y(
        N968) );
  OAI22X1TF U439 ( .A0(N188), .A1(N728), .B0(N794), .B1(N1047), .Y(N967) );
  OAI21X1TF U440 ( .A0(N738), .A1(N197), .B0(N1028), .Y(N5150) );
  AOI211X1TF U441 ( .A0(N1134), .A1(N284), .B0(N1027), .C0(N1026), .Y(N1028)
         );
  OAI22X1TF U442 ( .A0(N187), .A1(N720), .B0(N786), .B1(N1047), .Y(N1027) );
  OAI21X1TF U443 ( .A0(N747), .A1(N197), .B0(N987), .Y(N4730) );
  AOI211X1TF U444 ( .A0(N1134), .A1(IO_DATAOUTB[6]), .B0(N986), .C0(N985), .Y(
        N987) );
  OAI22X1TF U445 ( .A0(N811), .A1(N209), .B0(N779), .B1(N191), .Y(N985) );
  OAI22X1TF U446 ( .A0(N188), .A1(N729), .B0(N795), .B1(N1047), .Y(N986) );
  OAI21X1TF U447 ( .A0(N741), .A1(N197), .B0(N1037), .Y(N518) );
  AOI211X1TF U448 ( .A0(N200), .A1(IO_DATAOUTB[12]), .B0(N1036), .C0(N1035), 
        .Y(N1037) );
  OAI22X1TF U449 ( .A0(N805), .A1(N209), .B0(N773), .B1(N192), .Y(N1035) );
  OAI22X1TF U450 ( .A0(N1048), .A1(N723), .B0(N789), .B1(N1047), .Y(N1036) );
  OAI21X1TF U451 ( .A0(N742), .A1(N198), .B0(N1040), .Y(N519) );
  AOI211X1TF U452 ( .A0(N200), .A1(IO_DATAOUTB[11]), .B0(N1039), .C0(N1038), 
        .Y(N1040) );
  OAI22X1TF U453 ( .A0(N806), .A1(N209), .B0(N774), .B1(N192), .Y(N1038) );
  OAI22X1TF U454 ( .A0(N188), .A1(N724), .B0(N790), .B1(N1047), .Y(N1039) );
  OAI21X1TF U455 ( .A0(N750), .A1(N198), .B0(N993), .Y(N4770) );
  AOI211X1TF U456 ( .A0(N200), .A1(N995), .B0(N992), .C0(N991), .Y(N993) );
  OAI22X1TF U457 ( .A0(N814), .A1(N209), .B0(N782), .B1(N192), .Y(N991) );
  OAI22X1TF U458 ( .A0(N187), .A1(N732), .B0(N798), .B1(N205), .Y(N992) );
  OAI21X1TF U459 ( .A0(N739), .A1(N198), .B0(N1031), .Y(N5160) );
  AOI211X1TF U460 ( .A0(N200), .A1(N286), .B0(N1030), .C0(N1029), .Y(N1031) );
  OAI22X1TF U461 ( .A0(N188), .A1(N721), .B0(N787), .B1(N205), .Y(N1030) );
  OAI21X1TF U462 ( .A0(N745), .A1(N198), .B0(N1135), .Y(N522) );
  AOI211X1TF U463 ( .A0(N200), .A1(IO_DATAOUTB[8]), .B0(N1133), .C0(N1132), 
        .Y(N1135) );
  OAI22X1TF U464 ( .A0(N809), .A1(N209), .B0(N777), .B1(N192), .Y(N1132) );
  OAI22X1TF U465 ( .A0(N187), .A1(N727), .B0(N793), .B1(N205), .Y(N1133) );
  OAI21X1TF U466 ( .A0(N751), .A1(N198), .B0(N1000), .Y(N4800) );
  AOI211X1TF U467 ( .A0(N200), .A1(IO_DATAOUTB[2]), .B0(N999), .C0(N998), .Y(
        N1000) );
  OAI22X1TF U468 ( .A0(N815), .A1(N209), .B0(N783), .B1(N192), .Y(N998) );
  OAI22X1TF U469 ( .A0(N188), .A1(N733), .B0(N799), .B1(N205), .Y(N999) );
  OAI21X1TF U470 ( .A0(N748), .A1(N198), .B0(N984), .Y(N466) );
  AOI211X1TF U471 ( .A0(N200), .A1(IO_DATAOUTB[5]), .B0(N983), .C0(N982), .Y(
        N984) );
  OAI22X1TF U472 ( .A0(N812), .A1(N209), .B0(N780), .B1(N192), .Y(N982) );
  OAI22X1TF U473 ( .A0(N187), .A1(N730), .B0(N796), .B1(N205), .Y(N983) );
  OAI21X1TF U474 ( .A0(N752), .A1(N198), .B0(N1006), .Y(N4830) );
  AOI211X1TF U475 ( .A0(N200), .A1(N1008), .B0(N1005), .C0(N1004), .Y(N1006)
         );
  OAI22X1TF U476 ( .A0(N816), .A1(N209), .B0(N784), .B1(N192), .Y(N1004) );
  OAI22X1TF U477 ( .A0(N188), .A1(N734), .B0(N800), .B1(N205), .Y(N1005) );
  OAI21X1TF U478 ( .A0(N744), .A1(N198), .B0(N1046), .Y(N521) );
  AOI211X1TF U479 ( .A0(N200), .A1(IO_DATAOUTB[9]), .B0(N1045), .C0(N1044), 
        .Y(N1046) );
  OAI22X1TF U480 ( .A0(N808), .A1(N209), .B0(N776), .B1(N192), .Y(N1044) );
  OAI22X1TF U481 ( .A0(N188), .A1(N726), .B0(N792), .B1(N205), .Y(N1045) );
  AOI22X1TF U482 ( .A0(N190), .A1(N1143), .B0(N417), .B1(N1137), .Y(N530) );
  AOI22X1TF U483 ( .A0(N189), .A1(N1140), .B0(N403), .B1(N1137), .Y(N538) );
  AOI22X1TF U484 ( .A0(N190), .A1(N1141), .B0(N411), .B1(N1137), .Y(N536) );
  AOI22X1TF U485 ( .A0(N168), .A1(N1140), .B0(N263), .B1(N1142), .Y(N575) );
  INVX2TF U486 ( .A(I_DATAIN[7]), .Y(N1140) );
  AOI22X1TF U487 ( .A0(N168), .A1(N1141), .B0(N264), .B1(N1142), .Y(N577) );
  INVX2TF U488 ( .A(I_DATAIN[6]), .Y(N1141) );
  AOI22X1TF U489 ( .A0(N168), .A1(N1143), .B0(N53), .B1(N1142), .Y(N583) );
  INVX2TF U490 ( .A(I_DATAIN[3]), .Y(N1143) );
  AOI32X1TF U491 ( .A0(N572), .A1(N571), .A2(N203), .B0(N293), .B1(N571), .Y(
        N655) );
  AOI22X1TF U492 ( .A0(N570), .A1(N569), .B0(N576), .B1(D_ADDR[8]), .Y(N571)
         );
  INVX2TF U493 ( .A(N578), .Y(N569) );
  AOI22X1TF U494 ( .A0(N462), .A1(N4740), .B0(N756), .B1(N461), .Y(N1100) );
  AOI22X1TF U495 ( .A0(N444), .A1(N4680), .B0(N793), .B1(N443), .Y(N1121) );
  AOI22X1TF U496 ( .A0(N447), .A1(N4740), .B0(N772), .B1(N445), .Y(N1108) );
  AOI22X1TF U497 ( .A0(N485), .A1(N4720), .B0(N741), .B1(N4790), .Y(N1093) );
  AOI22X1TF U498 ( .A0(N485), .A1(N4680), .B0(N745), .B1(N4790), .Y(N1097) );
  AOI22X1TF U499 ( .A0(N485), .A1(N4700), .B0(N743), .B1(N4790), .Y(N1095) );
  AOI22X1TF U500 ( .A0(N485), .A1(N4710), .B0(N742), .B1(N4790), .Y(N1094) );
  AOI22X1TF U501 ( .A0(N485), .A1(N4690), .B0(N744), .B1(N4790), .Y(N1096) );
  AOI22X1TF U502 ( .A0(N485), .A1(N4740), .B0(N740), .B1(N4790), .Y(N1092) );
  AOI22X1TF U503 ( .A0(N442), .A1(N4690), .B0(N808), .B1(N441), .Y(N1128) );
  AOI22X1TF U504 ( .A0(N442), .A1(N4740), .B0(N804), .B1(N441), .Y(N1124) );
  AOI22X1TF U505 ( .A0(N442), .A1(N4720), .B0(N805), .B1(N441), .Y(N1125) );
  AOI22X1TF U506 ( .A0(N442), .A1(N4680), .B0(N809), .B1(N441), .Y(N1129) );
  AOI22X1TF U507 ( .A0(N442), .A1(N4710), .B0(N806), .B1(N441), .Y(N1126) );
  AOI22X1TF U508 ( .A0(N442), .A1(N4700), .B0(N807), .B1(N441), .Y(N1127) );
  AOI22X1TF U509 ( .A0(N447), .A1(N4820), .B0(N770), .B1(N445), .Y(N1106) );
  AOI22X1TF U510 ( .A0(N462), .A1(N4820), .B0(N754), .B1(N461), .Y(N1098) );
  AOI22X1TF U511 ( .A0(N462), .A1(N4760), .B0(N755), .B1(N461), .Y(N1099) );
  AOI22X1TF U512 ( .A0(N447), .A1(N4760), .B0(N771), .B1(N445), .Y(N1107) );
  AOI22X1TF U513 ( .A0(N499), .A1(N5050), .B0(N765), .B1(N498), .Y(N1061) );
  AOI22X1TF U514 ( .A0(N494), .A1(N5050), .B0(N797), .B1(N493), .Y(N1077) );
  AOI22X1TF U515 ( .A0(N494), .A1(N5030), .B0(N799), .B1(N493), .Y(N1079) );
  AOI22X1TF U516 ( .A0(N499), .A1(N5040), .B0(N766), .B1(N498), .Y(N1062) );
  AOI22X1TF U517 ( .A0(N499), .A1(N5060), .B0(N764), .B1(N498), .Y(N1060) );
  AOI22X1TF U518 ( .A0(N496), .A1(N5020), .B0(N784), .B1(N495), .Y(N1072) );
  AOI22X1TF U519 ( .A0(N496), .A1(N5030), .B0(N783), .B1(N495), .Y(N1071) );
  AOI22X1TF U520 ( .A0(N496), .A1(N5060), .B0(N780), .B1(N495), .Y(N1068) );
  AOI22X1TF U521 ( .A0(N494), .A1(N5010), .B0(N801), .B1(N493), .Y(N1081) );
  INVX2TF U522 ( .A(N494), .Y(N493) );
  AOI22X1TF U523 ( .A0(N485), .A1(N4820), .B0(N738), .B1(N4790), .Y(N1090) );
  AOI22X1TF U524 ( .A0(N442), .A1(N4820), .B0(N802), .B1(N441), .Y(N1122) );
  AOI22X1TF U525 ( .A0(N485), .A1(N4760), .B0(N739), .B1(N4790), .Y(N1091) );
  NAND4X2TF U526 ( .A(N4670), .B(N265), .C(N696), .D(N697), .Y(N4790) );
  AOI22X1TF U527 ( .A0(N442), .A1(N4760), .B0(N803), .B1(N441), .Y(N1123) );
  INVX2TF U528 ( .A(N488), .Y(N440) );
  NAND2X2TF U529 ( .A(N4670), .B(N964), .Y(N441) );
  AOI22X1TF U530 ( .A0(N5100), .A1(N5090), .B0(N746), .B1(N5080), .Y(N1050) );
  AOI22X1TF U531 ( .A0(N491), .A1(N5090), .B0(N810), .B1(N490), .Y(N1082) );
  AOI22X1TF U532 ( .A0(N5100), .A1(N5070), .B0(N747), .B1(N5080), .Y(N1051) );
  AOI22X1TF U533 ( .A0(N5100), .A1(N5050), .B0(N749), .B1(N5080), .Y(N1053) );
  AOI22X1TF U534 ( .A0(N5100), .A1(N5030), .B0(N751), .B1(N5080), .Y(N1055) );
  AOI22X1TF U535 ( .A0(N5100), .A1(N5020), .B0(N752), .B1(N5080), .Y(N1056) );
  AOI22X1TF U536 ( .A0(N5100), .A1(N5040), .B0(N750), .B1(N5080), .Y(N1054) );
  AOI22X1TF U537 ( .A0(N5100), .A1(N5060), .B0(N748), .B1(N5080), .Y(N1052) );
  AOI22X1TF U538 ( .A0(N5100), .A1(N5010), .B0(N753), .B1(N5080), .Y(N1057) );
  NAND4X2TF U539 ( .A(N500), .B(N265), .C(N696), .D(N697), .Y(N5080) );
  AOI22X1TF U540 ( .A0(N491), .A1(N5070), .B0(N811), .B1(N490), .Y(N1083) );
  AOI22X1TF U541 ( .A0(N491), .A1(N5050), .B0(N813), .B1(N490), .Y(N1085) );
  AOI22X1TF U542 ( .A0(N491), .A1(N5030), .B0(N815), .B1(N490), .Y(N1087) );
  AOI22X1TF U543 ( .A0(N491), .A1(N5020), .B0(N816), .B1(N490), .Y(N1088) );
  AOI22X1TF U544 ( .A0(N491), .A1(N5060), .B0(N812), .B1(N490), .Y(N1084) );
  AOI22X1TF U545 ( .A0(N491), .A1(N5040), .B0(N814), .B1(N490), .Y(N1086) );
  AOI22X1TF U546 ( .A0(N491), .A1(N5010), .B0(N817), .B1(N490), .Y(N1089) );
  NAND2X2TF U547 ( .A(N500), .B(N964), .Y(N490) );
  AOI32X4TF U548 ( .A0(N580), .A1(N487), .A2(N423), .B0(N438), .B1(N487), .Y(
        N488) );
  OAI211X1TF U549 ( .A0(N429), .A1(N937), .B0(N971), .C0(N437), .Y(N438) );
  OAI211X1TF U550 ( .A0(N1178), .A1(N1225), .B0(N1158), .C0(N1157), .Y(N601)
         );
  AOI22X1TF U551 ( .A0(IO_DATAINA[8]), .A1(N298), .B0(N395), .B1(N1156), .Y(
        N1157) );
  OAI211X1TF U552 ( .A0(N399), .A1(N1225), .B0(N1186), .C0(N1185), .Y(N617) );
  AOI22X1TF U553 ( .A0(IO_DATAINA[3]), .A1(N397), .B0(N395), .B1(N1184), .Y(
        N1185) );
  AOI22X1TF U554 ( .A0(IO_DATAINB[3]), .A1(N199), .B0(D_ADDR[4]), .B1(N1238), 
        .Y(N1186) );
  OAI211X1TF U555 ( .A0(N1171), .A1(N1225), .B0(N1170), .C0(N1169), .Y(N609)
         );
  AOI22X1TF U556 ( .A0(IO_DATAINA[4]), .A1(N298), .B0(N395), .B1(N1183), .Y(
        N1169) );
  INVX2TF U557 ( .A(N399), .Y(N1183) );
  AOI22X1TF U558 ( .A0(IO_DATAINB[4]), .A1(N398), .B0(D_ADDR[5]), .B1(N296), 
        .Y(N1170) );
  OAI211X1TF U559 ( .A0(N1165), .A1(N1224), .B0(N1145), .C0(N1144), .Y(N593)
         );
  AOI22X1TF U560 ( .A0(IO_DATAINA[7]), .A1(N298), .B0(N396), .B1(N1156), .Y(
        N1144) );
  AOI22X1TF U561 ( .A0(IO_DATAINB[7]), .A1(N199), .B0(D_ADDR[8]), .B1(N1238), 
        .Y(N1145) );
  OAI31X1TF U562 ( .A0(I_ADDR[2]), .A1(N292), .A2(N203), .B0(N568), .Y(N656)
         );
  AOI22X1TF U563 ( .A0(I_ADDR[2]), .A1(N567), .B0(N576), .B1(D_ADDR[2]), .Y(
        N568) );
  OAI21X1TF U564 ( .A0(I_ADDR[1]), .A1(N578), .B0(N572), .Y(N567) );
  OAI31X1TF U565 ( .A0(I_ADDR[4]), .A1(N566), .A2(N203), .B0(N565), .Y(N658)
         );
  AOI22X1TF U566 ( .A0(I_ADDR[4]), .A1(N564), .B0(N576), .B1(D_ADDR[4]), .Y(
        N565) );
  OAI21X1TF U567 ( .A0(N563), .A1(N578), .B0(N572), .Y(N564) );
  OAI31X1TF U568 ( .A0(I_ADDR[6]), .A1(N561), .A2(N203), .B0(N560), .Y(N660)
         );
  AOI22X1TF U569 ( .A0(I_ADDR[6]), .A1(N559), .B0(N576), .B1(D_ADDR[6]), .Y(
        N560) );
  OAI211X1TF U570 ( .A0(N401), .A1(N1225), .B0(N1139), .C0(N1138), .Y(N573) );
  AOI22X1TF U571 ( .A0(IO_DATAINA[10]), .A1(N298), .B0(N395), .B1(N1175), .Y(
        N1138) );
  OAI211X1TF U572 ( .A0(N1178), .A1(N1224), .B0(N1177), .C0(N1176), .Y(N613)
         );
  AOI22X1TF U573 ( .A0(IO_DATAINA[9]), .A1(N298), .B0(N396), .B1(N1175), .Y(
        N1176) );
  OAI211X1TF U574 ( .A0(N1165), .A1(N1225), .B0(N1164), .C0(N1163), .Y(N605)
         );
  AOI22X1TF U575 ( .A0(IO_DATAINB[6]), .A1(N199), .B0(D_ADDR[7]), .B1(N1238), 
        .Y(N1164) );
  OAI211X1TF U576 ( .A0(N1171), .A1(N1224), .B0(N973), .C0(N972), .Y(N463) );
  AOI22X1TF U577 ( .A0(IO_DATAINB[5]), .A1(N398), .B0(D_ADDR[6]), .B1(N296), 
        .Y(N973) );
  OAI211X1TF U578 ( .A0(N401), .A1(N1224), .B0(N1198), .C0(N1197), .Y(N625) );
  AOI22X1TF U579 ( .A0(IO_DATAINA[11]), .A1(N397), .B0(N396), .B1(N1196), .Y(
        N1197) );
  OAI211X1TF U580 ( .A0(N400), .A1(N1225), .B0(N1191), .C0(N1190), .Y(N621) );
  AOI22X1TF U581 ( .A0(IO_DATAINA[12]), .A1(N397), .B0(N395), .B1(N1196), .Y(
        N1190) );
  OAI211X1TF U582 ( .A0(N1152), .A1(N1224), .B0(N1151), .C0(N1150), .Y(N597)
         );
  AOI22X1TF U583 ( .A0(IO_DATAINA[2]), .A1(N298), .B0(N396), .B1(N1184), .Y(
        N1150) );
  AOI22X1TF U584 ( .A0(IO_DATAINB[2]), .A1(N199), .B0(D_ADDR[3]), .B1(N1238), 
        .Y(N1151) );
  INVX2TF U585 ( .A(N1207), .Y(N1152) );
  OAI211X1TF U586 ( .A0(N177), .A1(N816), .B0(N1010), .C0(N1009), .Y(N484) );
  AOI21X1TF U587 ( .A0(N1008), .A1(N175), .B0(N1007), .Y(N1009) );
  INVX2TF U588 ( .A(N768), .Y(N1008) );
  AOI22X1TF U589 ( .A0(IO_DATAOUTA[1]), .A1(N1015), .B0(N1016), .B1(
        IO_OFFSET[1]), .Y(N1010) );
  OAI211X1TF U590 ( .A0(N177), .A1(N815), .B0(N1003), .C0(N1002), .Y(N4810) );
  AOI21X1TF U591 ( .A0(IO_DATAOUTB[2]), .A1(N175), .B0(N1001), .Y(N1002) );
  AOI22X1TF U592 ( .A0(IO_DATAOUTA[2]), .A1(N1015), .B0(N1016), .B1(
        IO_OFFSET[2]), .Y(N1003) );
  OAI211X1TF U593 ( .A0(N177), .A1(N810), .B0(N959), .C0(N958), .Y(N459) );
  AOI21X1TF U594 ( .A0(IO_DATAOUTB[7]), .A1(N175), .B0(N957), .Y(N958) );
  AOI22X1TF U595 ( .A0(IO_DATAOUTA[7]), .A1(N1015), .B0(N1016), .B1(
        IO_OFFSET[7]), .Y(N959) );
  OAI211X1TF U596 ( .A0(N177), .A1(N814), .B0(N997), .C0(N996), .Y(N4780) );
  AOI21X1TF U597 ( .A0(N995), .A1(N175), .B0(N994), .Y(N996) );
  INVX2TF U598 ( .A(N766), .Y(N995) );
  AOI22X1TF U599 ( .A0(IO_DATAOUTA[3]), .A1(N1015), .B0(N1016), .B1(
        IO_OFFSET[3]), .Y(N997) );
  OAI211X1TF U600 ( .A0(N177), .A1(N812), .B0(N981), .C0(N980), .Y(N465) );
  AOI21X1TF U601 ( .A0(IO_DATAOUTB[5]), .A1(N175), .B0(N979), .Y(N980) );
  AOI22X1TF U602 ( .A0(IO_DATAOUTA[5]), .A1(N1015), .B0(N1016), .B1(
        IO_OFFSET[5]), .Y(N981) );
  OAI21X1TF U603 ( .A0(N578), .A1(N558), .B0(N572), .Y(N559) );
  INVX2TF U604 ( .A(N574), .Y(N572) );
  NOR2X2TF U605 ( .A(N553), .B(N552), .Y(N576) );
  AOI32X1TF U606 ( .A0(N550), .A1(N939), .A2(CF), .B0(N549), .B1(N939), .Y(
        N552) );
  OAI211X1TF U607 ( .A0(CF), .A1(N894), .B0(N548), .C0(N547), .Y(N549) );
  OAI21X1TF U608 ( .A0(N169), .A1(NF), .B0(CODE_TYPE[2]), .Y(N546) );
  AOI32X1TF U609 ( .A0(N169), .A1(ZF), .A2(N55), .B0(N940), .B1(N290), .Y(N548) );
  INVX2TF U610 ( .A(N566), .Y(N563) );
  AOI21X1TF U611 ( .A0(N298), .A1(IO_DATAINA[13]), .B0(N1202), .Y(N1203) );
  OAI22X1TF U612 ( .A0(N400), .A1(N1224), .B0(N410), .B1(N414), .Y(N1202) );
  OAI211X1TF U613 ( .A0(N402), .A1(N1224), .B0(N1205), .C0(N1204), .Y(N1206)
         );
  AOI22X1TF U614 ( .A0(N298), .A1(IO_DATAINA[1]), .B0(N394), .B1(IO_STATUS[1]), 
        .Y(N1204) );
  AOI22X1TF U615 ( .A0(IO_DATAINB[1]), .A1(N398), .B0(D_ADDR[2]), .B1(N296), 
        .Y(N1205) );
  OAI21X1TF U616 ( .A0(N177), .A1(N803), .B0(N1214), .Y(N634) );
  AOI211X1TF U617 ( .A0(N286), .A1(N174), .B0(N1212), .C0(N1211), .Y(N1214) );
  OAI21X1TF U618 ( .A0(N177), .A1(N807), .B0(N1025), .Y(N5140) );
  AOI211X1TF U619 ( .A0(IO_DATAOUTB[10]), .A1(N174), .B0(N1024), .C0(N1023), 
        .Y(N1025) );
  OAI22X1TF U620 ( .A0(N775), .A1(N1210), .B0(N1209), .B1(N743), .Y(N1023) );
  OAI21X1TF U621 ( .A0(N178), .A1(N809), .B0(N1155), .Y(N598) );
  AOI211X1TF U622 ( .A0(IO_DATAOUTB[8]), .A1(N174), .B0(N1154), .C0(N1153), 
        .Y(N1155) );
  OAI22X1TF U623 ( .A0(N777), .A1(N1210), .B0(N1209), .B1(N745), .Y(N1153) );
  OAI21X1TF U624 ( .A0(N178), .A1(N805), .B0(N1189), .Y(N618) );
  AOI211X1TF U625 ( .A0(IO_DATAOUTB[12]), .A1(N174), .B0(N1188), .C0(N1187), 
        .Y(N1189) );
  OAI22X1TF U626 ( .A0(N773), .A1(N1210), .B0(N1209), .B1(N741), .Y(N1187) );
  OAI21X1TF U627 ( .A0(N178), .A1(N806), .B0(N1022), .Y(N5130) );
  AOI211X1TF U628 ( .A0(IO_DATAOUTB[11]), .A1(N174), .B0(N1021), .C0(N1020), 
        .Y(N1022) );
  OAI22X1TF U629 ( .A0(N774), .A1(N1210), .B0(N1209), .B1(N742), .Y(N1020) );
  OAI21X1TF U630 ( .A0(N178), .A1(N804), .B0(N1201), .Y(N626) );
  AOI211X1TF U631 ( .A0(N285), .A1(N174), .B0(N1200), .C0(N1199), .Y(N1201) );
  OAI21X1TF U632 ( .A0(N178), .A1(N808), .B0(N1174), .Y(N610) );
  AOI211X1TF U633 ( .A0(IO_DATAOUTB[9]), .A1(N174), .B0(N1173), .C0(N1172), 
        .Y(N1174) );
  OAI22X1TF U634 ( .A0(N776), .A1(N1210), .B0(N1209), .B1(N744), .Y(N1172) );
  OAI21X1TF U635 ( .A0(N178), .A1(N802), .B0(N1019), .Y(N5120) );
  AOI211X1TF U636 ( .A0(N284), .A1(N175), .B0(N1018), .C0(N1017), .Y(N1019) );
  OAI21X1TF U637 ( .A0(N178), .A1(N813), .B0(N1168), .Y(N606) );
  AOI211X1TF U638 ( .A0(IO_DATAOUTB[4]), .A1(N174), .B0(N1167), .C0(N1166), 
        .Y(N1168) );
  OAI22X1TF U639 ( .A0(N781), .A1(N1210), .B0(N1209), .B1(N749), .Y(N1166) );
  OAI21X1TF U640 ( .A0(N178), .A1(N811), .B0(N1161), .Y(N602) );
  AOI211X1TF U641 ( .A0(IO_DATAOUTB[6]), .A1(N175), .B0(N1160), .C0(N1159), 
        .Y(N1161) );
  OAI22X1TF U642 ( .A0(N779), .A1(N1210), .B0(N1209), .B1(N747), .Y(N1159) );
  OAI22X2TF U643 ( .A0(N695), .A1(N948), .B0(N411), .B1(N950), .Y(N1016) );
  INVX2TF U644 ( .A(N1015), .Y(N1210) );
  OAI2BB2X2TF U645 ( .B0(N413), .B1(N946), .A0N(N965), .A1N(N952), .Y(N1015)
         );
  OAI31X1TF U646 ( .A0(N955), .A1(N954), .A2(N953), .B0(N961), .Y(N956) );
  NOR2X1TF U647 ( .A(N412), .B(N950), .Y(N951) );
  INVX2TF U648 ( .A(N950), .Y(N947) );
  AND2X2TF U649 ( .A(N964), .B(N952), .Y(N944) );
  AOI22X1TF U650 ( .A0(CODE_TYPE[3]), .A1(N940), .B0(N939), .B1(N938), .Y(N942) );
  INVX2TF U651 ( .A(N893), .Y(N939) );
  AOI22X1TF U652 ( .A0(IO_DATAINA[14]), .A1(N397), .B0(N396), .B1(N1237), .Y(
        N1216) );
  AOI22X1TF U653 ( .A0(N395), .A1(N1223), .B0(REG_C[14]), .B1(N1238), .Y(N1217) );
  AOI22X1TF U654 ( .A0(N397), .A1(IO_DATAINA[15]), .B0(REG_C[15]), .B1(N296), 
        .Y(N392) );
  OAI22X1TF U655 ( .A0(N889), .A1(N888), .B0(N290), .B1(N409), .Y(N450) );
  OR4X2TF U656 ( .A(N859), .B(N346), .C(N858), .D(N345), .Y(N1156) );
  AOI22X1TF U657 ( .A0(N850), .A1(N851), .B0(N405), .B1(N860), .Y(N344) );
  OAI21X1TF U658 ( .A0(N857), .A1(N856), .B0(N855), .Y(N858) );
  AOI22X1TF U659 ( .A0(N406), .A1(N854), .B0(N1630), .B1(N853), .Y(N855) );
  AOI21X1TF U660 ( .A0(N204), .A1(N343), .B0(N215), .Y(N346) );
  AOI22X1TF U661 ( .A0(N420), .A1(N272), .B0(N295), .B1(REG_A[7]), .Y(N343) );
  AOI21X1TF U662 ( .A0(N303), .A1(N215), .B0(N876), .Y(N852) );
  OAI211X1TF U663 ( .A0(N703), .A1(N848), .B0(N702), .C0(N701), .Y(N1207) );
  AOI32X1TF U664 ( .A0(N302), .A1(REG_A[1]), .A2(N210), .B0(N823), .B1(
        REG_A[1]), .Y(N701) );
  OAI31X1TF U665 ( .A0(N834), .A1(REG_B[3]), .A2(N885), .B0(N318), .Y(N319) );
  AOI31X1TF U666 ( .A0(N692), .A1(N691), .A2(N690), .B0(N827), .Y(N699) );
  AND2X2TF U667 ( .A(N719), .B(N329), .Y(N399) );
  AOI21X1TF U668 ( .A0(N470), .A1(N159), .B0(N326), .Y(N327) );
  OAI211X1TF U669 ( .A0(N279), .A1(N166), .B0(N708), .C0(N707), .Y(N709) );
  AOI22X1TF U670 ( .A0(N851), .A1(N853), .B0(N714), .B1(N850), .Y(N736) );
  AOI221X1TF U671 ( .A0(N273), .A1(N302), .B0(REG_A[3]), .B1(N295), .C0(N716), 
        .Y(N717) );
  OAI31X1TF U672 ( .A0(N848), .A1(N57), .A2(N857), .B0(N838), .Y(N716) );
  OAI21X1TF U673 ( .A0(REG_B[3]), .A1(N879), .B0(N715), .Y(N718) );
  OR2X2TF U674 ( .A(N826), .B(N335), .Y(N1184) );
  OAI21X1TF U675 ( .A0(N820), .A1(N211), .B0(N334), .Y(N335) );
  AOI211X1TF U676 ( .A0(REG_A[4]), .A1(N183), .B0(N818), .C0(N737), .Y(N828)
         );
  OAI22X1TF U677 ( .A0(N825), .A1(N271), .B0(N824), .B1(N57), .Y(N826) );
  AOI221X1TF U678 ( .A0(N302), .A1(N271), .B0(N421), .B1(REG_A[2]), .C0(N881), 
        .Y(N824) );
  AOI21X1TF U679 ( .A0(N302), .A1(N57), .B0(N823), .Y(N825) );
  INVX2TF U680 ( .A(N715), .Y(N823) );
  AOI21X1TF U681 ( .A0(N476), .A1(N180), .B0(N341), .Y(N342) );
  AOI22X1TF U682 ( .A0(N829), .A1(N406), .B0(N405), .B1(N837), .Y(N338) );
  INVX2TF U683 ( .A(N835), .Y(N339) );
  OAI31X1TF U684 ( .A0(N211), .A1(N885), .A2(N834), .B0(N833), .Y(N835) );
  AOI22X1TF U685 ( .A0(N1630), .A1(N832), .B0(N851), .B1(N831), .Y(N833) );
  INVX2TF U686 ( .A(N688), .Y(N831) );
  AOI21X1TF U687 ( .A0(N302), .A1(N217), .B0(N876), .Y(N830) );
  OAI211X1TF U688 ( .A0(N278), .A1(N166), .B0(N705), .C0(N704), .Y(N850) );
  AOI21X1TF U689 ( .A0(N481), .A1(N180), .B0(N320), .Y(N321) );
  OAI21X1TF U690 ( .A0(N886), .A1(N885), .B0(N884), .Y(N320) );
  OAI32X1TF U691 ( .A0(N883), .A1(N882), .A2(N881), .B0(REG_B[14]), .B1(N883), 
        .Y(N884) );
  AOI22X1TF U692 ( .A0(REG_A[14]), .A1(N880), .B0(N879), .B1(N278), .Y(N882)
         );
  OAI31X1TF U693 ( .A0(REG_B[2]), .A1(REG_B[3]), .A2(N878), .B0(N877), .Y(N883) );
  AOI32X1TF U694 ( .A0(N302), .A1(REG_A[14]), .A2(N222), .B0(N876), .B1(
        REG_A[14]), .Y(N877) );
  INVX2TF U695 ( .A(N875), .Y(N878) );
  AOI211X1TF U696 ( .A0(N428), .A1(N873), .B0(N872), .C0(N871), .Y(N886) );
  AOI31X1TF U697 ( .A0(N866), .A1(N865), .A2(N864), .B0(N863), .Y(N872) );
  INVX2TF U698 ( .A(N861), .Y(N873) );
  AOI211X1TF U699 ( .A0(N851), .A1(N832), .B0(N640), .C0(N639), .Y(N1162) );
  OAI211X1TF U700 ( .A0(N317), .A1(N213), .B0(N636), .C0(N316), .Y(N639) );
  AOI22X1TF U701 ( .A0(N506), .A1(N874), .B0(N472), .B1(N159), .Y(N316) );
  AOI22X1TF U702 ( .A0(REG_A[5]), .A1(N635), .B0(N1630), .B1(N689), .Y(N636)
         );
  AOI211X1TF U703 ( .A0(N303), .A1(N282), .B0(N881), .C0(N315), .Y(N317) );
  NOR2X1TF U704 ( .A(N880), .B(N282), .Y(N315) );
  OAI22X1TF U705 ( .A0(N688), .A1(N856), .B0(N682), .B1(N628), .Y(N640) );
  NOR2X1TF U706 ( .A(N848), .B(N652), .Y(N875) );
  INVX2TF U707 ( .A(N822), .Y(N870) );
  INVX2TF U708 ( .A(N856), .Y(N714) );
  NOR2X2TF U709 ( .A(N595), .B(N848), .Y(N851) );
  OAI21X1TF U710 ( .A0(N748), .A1(N196), .B0(N978), .Y(N464) );
  NOR3X1TF U711 ( .A(N977), .B(N976), .C(N975), .Y(N978) );
  OAI22X1TF U712 ( .A0(N796), .A1(N182), .B0(N213), .B1(N1236), .Y(N975) );
  OAI22X1TF U713 ( .A0(N413), .A1(N974), .B0(N764), .B1(N1227), .Y(N977) );
  OAI21X1TF U714 ( .A0(N749), .A1(N196), .B0(N921), .Y(N455) );
  NOR3X1TF U715 ( .A(N920), .B(N919), .C(N918), .Y(N921) );
  OAI22X1TF U716 ( .A0(N797), .A1(N182), .B0(N212), .B1(N1236), .Y(N918) );
  OAI22X1TF U717 ( .A0(N412), .A1(N974), .B0(N765), .B1(N1227), .Y(N920) );
  OAI21X1TF U718 ( .A0(N750), .A1(N196), .B0(N1182), .Y(N614) );
  NOR3X1TF U719 ( .A(N1181), .B(N1180), .C(N1179), .Y(N1182) );
  OAI22X1TF U720 ( .A0(N798), .A1(N182), .B0(N211), .B1(N1236), .Y(N1179) );
  OAI22X1TF U721 ( .A0(N766), .A1(N1227), .B0(N417), .B1(N1218), .Y(N1181) );
  OAI21X1TF U722 ( .A0(N751), .A1(N196), .B0(N1149), .Y(N594) );
  NOR3X1TF U723 ( .A(N1148), .B(N1147), .C(N1146), .Y(N1149) );
  OAI22X1TF U724 ( .A0(N799), .A1(N182), .B0(N57), .B1(N1236), .Y(N1146) );
  OAI22X1TF U725 ( .A0(N767), .A1(N1227), .B0(N269), .B1(N1218), .Y(N1148) );
  OAI21X1TF U726 ( .A0(N747), .A1(N196), .B0(N925), .Y(N456) );
  NOR3X1TF U727 ( .A(N924), .B(N923), .C(N922), .Y(N925) );
  OAI22X1TF U728 ( .A0(N795), .A1(N182), .B0(N214), .B1(N1236), .Y(N922) );
  OAI22X1TF U729 ( .A0(N811), .A1(N171), .B0(N779), .B1(N194), .Y(N923) );
  OAI22X1TF U730 ( .A0(N411), .A1(N974), .B0(N763), .B1(N1227), .Y(N924) );
  OAI21X1TF U731 ( .A0(N746), .A1(N196), .B0(N933), .Y(N458) );
  NOR3X1TF U732 ( .A(N932), .B(N931), .C(N930), .Y(N933) );
  OAI22X1TF U733 ( .A0(N794), .A1(N182), .B0(N215), .B1(N1236), .Y(N930) );
  OAI22X1TF U734 ( .A0(N810), .A1(N171), .B0(N778), .B1(N194), .Y(N931) );
  OAI22X1TF U735 ( .A0(N762), .A1(N201), .B0(N403), .B1(N974), .Y(N932) );
  OAI21X1TF U736 ( .A0(N753), .A1(N196), .B0(N1222), .Y(N638) );
  NOR3X1TF U737 ( .A(N1221), .B(N1220), .C(N1219), .Y(N1222) );
  OAI22X1TF U738 ( .A0(N801), .A1(N182), .B0(N54), .B1(N1236), .Y(N1219) );
  OAI22X1TF U739 ( .A0(N817), .A1(N171), .B0(N785), .B1(N194), .Y(N1220) );
  OAI22X1TF U740 ( .A0(N769), .A1(N201), .B0(N259), .B1(N1218), .Y(N1221) );
  OAI21X1TF U741 ( .A0(N219), .A1(N206), .B0(N1195), .Y(N622) );
  NOR3X1TF U742 ( .A(N1194), .B(N1193), .C(N1192), .Y(N1195) );
  OAI22X1TF U743 ( .A0(N806), .A1(N171), .B0(N774), .B1(N193), .Y(N1193) );
  OAI22X1TF U744 ( .A0(N758), .A1(N201), .B0(N417), .B1(N1226), .Y(N1194) );
  OAI21X1TF U745 ( .A0(N221), .A1(N206), .B0(N908), .Y(N452) );
  NOR3X1TF U746 ( .A(N907), .B(N906), .C(N905), .Y(N908) );
  OAI22X1TF U747 ( .A0(N413), .A1(N1226), .B0(N756), .B1(N1227), .Y(N907) );
  OAI21X1TF U748 ( .A0(N217), .A1(N206), .B0(N916), .Y(N454) );
  NOR3X1TF U749 ( .A(N915), .B(N914), .C(N913), .Y(N916) );
  OAI22X1TF U750 ( .A0(N808), .A1(N170), .B0(N776), .B1(N194), .Y(N914) );
  OAI22X1TF U751 ( .A0(N760), .A1(N201), .B0(N261), .B1(N1226), .Y(N915) );
  OAI21X1TF U752 ( .A0(N216), .A1(N206), .B0(N929), .Y(N457) );
  NOR3X1TF U753 ( .A(N928), .B(N927), .C(N926), .Y(N929) );
  OAI22X1TF U754 ( .A0(N809), .A1(N170), .B0(N777), .B1(N194), .Y(N927) );
  OAI22X1TF U755 ( .A0(N761), .A1(N201), .B0(N259), .B1(N1226), .Y(N928) );
  OAI21X1TF U756 ( .A0(N223), .A1(N206), .B0(N1235), .Y(N642) );
  NOR3X1TF U757 ( .A(N1234), .B(N1233), .C(N1232), .Y(N1235) );
  OAI22X1TF U758 ( .A0(N754), .A1(N201), .B0(N403), .B1(N1226), .Y(N1234) );
  OAI21X1TF U759 ( .A0(N220), .A1(N206), .B0(N912), .Y(N453) );
  NOR3X1TF U760 ( .A(N911), .B(N910), .C(N909), .Y(N912) );
  OAI22X1TF U761 ( .A0(N805), .A1(N171), .B0(N773), .B1(N194), .Y(N910) );
  OAI22X1TF U762 ( .A0(N412), .A1(N1226), .B0(N757), .B1(N1227), .Y(N911) );
  OAI21X1TF U763 ( .A0(N222), .A1(N206), .B0(N904), .Y(N451) );
  NOR3X1TF U764 ( .A(N903), .B(N902), .C(N901), .Y(N904) );
  OAI22X1TF U765 ( .A0(N411), .A1(N1226), .B0(N755), .B1(N1227), .Y(N903) );
  NOR2X1TF U766 ( .A(OPER3_R3[1]), .B(N899), .Y(N900) );
  NOR2X1TF U767 ( .A(OPER3_R3[0]), .B(N899), .Y(N897) );
  INVX2TF U768 ( .A(N898), .Y(N899) );
  NAND2X2TF U769 ( .A(N891), .B(N961), .Y(N1226) );
  AOI21X1TF U770 ( .A0(N960), .A1(N943), .B0(N970), .Y(N891) );
  OAI211X1TF U771 ( .A0(CODE_TYPE[3]), .A1(N422), .B0(N961), .C0(N263), .Y(
        N896) );
  AOI21X1TF U772 ( .A0(IO_DATAINA[0]), .A1(N397), .B0(N388), .Y(N389) );
  OAI211X1TF U773 ( .A0(N402), .A1(N1225), .B0(N387), .C0(N386), .Y(N388) );
  AND2X2TF U774 ( .A(N383), .B(N422), .Y(N398) );
  AOI22X1TF U775 ( .A0(N394), .A1(IO_STATUS[0]), .B0(D_ADDR[1]), .B1(N296), 
        .Y(N387) );
  AOI21X1TF U776 ( .A0(N263), .A1(N169), .B0(N971), .Y(N381) );
  AOI211X1TF U777 ( .A0(\SUB_X_276_4_B[0] ), .A1(N375), .B0(N374), .C0(N373), 
        .Y(N402) );
  OAI211X1TF U778 ( .A0(N848), .A1(N849), .B0(N847), .C0(N372), .Y(N373) );
  AOI22X1TF U779 ( .A0(N159), .A1(N467), .B0(N501), .B1(N874), .Y(N372) );
  OAI31X1TF U780 ( .A0(N846), .A1(N845), .A2(N844), .B0(N162), .Y(N847) );
  NOR2X1TF U781 ( .A(N843), .B(N271), .Y(N844) );
  NOR2X1TF U782 ( .A(N842), .B(N59), .Y(N846) );
  INVX2TF U783 ( .A(N408), .Y(N848) );
  NOR2X1TF U784 ( .A(N370), .B(N1014), .Y(N374) );
  AOI21X1TF U785 ( .A0(N420), .A1(N54), .B0(N369), .Y(N370) );
  OAI211X1TF U786 ( .A0(REG_A[0]), .A1(N879), .B0(N838), .C0(N368), .Y(N375)
         );
  AOI21X1TF U787 ( .A0(N511), .A1(N874), .B0(N367), .Y(N401) );
  OAI211X1TF U788 ( .A0(N218), .A1(N366), .B0(N365), .C0(N665), .Y(N367) );
  AOI211X1TF U789 ( .A0(N406), .A1(N868), .B0(N664), .C0(N663), .Y(N665) );
  OAI22X1TF U790 ( .A0(N822), .A1(N662), .B0(REG_B[3]), .B1(N820), .Y(N663) );
  OAI211X1TF U791 ( .A0(N277), .A1(N166), .B0(N616), .C0(N667), .Y(N650) );
  AOI22X1TF U792 ( .A0(REG_A[10]), .A1(N347), .B0(N183), .B1(REG_A[12]), .Y(
        N616) );
  OAI22X1TF U793 ( .A0(N843), .A1(N1014), .B0(N842), .B1(N59), .Y(N611) );
  OAI22X1TF U794 ( .A0(N648), .A1(N283), .B0(N861), .B1(N821), .Y(N664) );
  NOR4X1TF U795 ( .A(N647), .B(N646), .C(N644), .D(N643), .Y(N861) );
  NOR2X1TF U796 ( .A(N283), .B(N675), .Y(N643) );
  NOR2X1TF U797 ( .A(N842), .B(N266), .Y(N644) );
  NOR2X1TF U798 ( .A(N843), .B(N274), .Y(N646) );
  NOR2X1TF U799 ( .A(N1650), .B(N272), .Y(N647) );
  AOI21X1TF U800 ( .A0(N218), .A1(N303), .B0(N876), .Y(N648) );
  NOR2X1TF U801 ( .A(N166), .B(N273), .Y(N845) );
  AOI211X1TF U802 ( .A0(N420), .A1(N283), .B0(N881), .C0(N364), .Y(N366) );
  NOR2X1TF U803 ( .A(N880), .B(N283), .Y(N364) );
  INVX2TF U804 ( .A(N295), .Y(N880) );
  OAI211X1TF U805 ( .A0(N673), .A1(N885), .B0(N362), .C0(N361), .Y(N363) );
  AOI21X1TF U806 ( .A0(N839), .A1(N1630), .B0(N360), .Y(N361) );
  OAI21X1TF U807 ( .A0(N359), .A1(N276), .B0(N358), .Y(N360) );
  AOI221X1TF U808 ( .A0(N302), .A1(N276), .B0(N295), .B1(REG_A[12]), .C0(N881), 
        .Y(N672) );
  OAI211X1TF U809 ( .A0(N266), .A1(N166), .B0(N667), .C0(N666), .Y(N668) );
  AOI21X1TF U810 ( .A0(N420), .A1(N220), .B0(N683), .Y(N359) );
  OAI211X1TF U811 ( .A0(N276), .A1(N675), .B0(N865), .C0(N592), .Y(N839) );
  AOI22X1TF U812 ( .A0(N56), .A1(REG_A[15]), .B0(N183), .B1(REG_A[14]), .Y(
        N592) );
  INVX2TF U813 ( .A(N407), .Y(N885) );
  NOR2X1TF U814 ( .A(N1650), .B(N282), .Y(N737) );
  NOR2X1TF U815 ( .A(N675), .B(N1014), .Y(N670) );
  OAI211X1TF U816 ( .A0(N59), .A1(N166), .B0(N599), .C0(N596), .Y(N671) );
  INVX2TF U817 ( .A(N818), .Y(N596) );
  NOR2X1TF U818 ( .A(N842), .B(N273), .Y(N818) );
  AOI211X1TF U819 ( .A0(N480), .A1(N180), .B0(N686), .C0(N324), .Y(N325) );
  AOI22X1TF U820 ( .A0(N405), .A1(N322), .B0(N837), .B1(N406), .Y(N323) );
  OAI211X1TF U821 ( .A0(N843), .A1(N287), .B0(N704), .C0(N712), .Y(N322) );
  OAI22X1TF U822 ( .A0(N682), .A1(N681), .B0(N688), .B1(N827), .Y(N687) );
  OAI22X1TF U823 ( .A0(N843), .A1(N267), .B0(N842), .B1(N278), .Y(N624) );
  AOI22X1TF U824 ( .A0(REG_B[2]), .A1(N694), .B0(N829), .B1(N57), .Y(N682) );
  OAI211X1TF U825 ( .A0(N271), .A1(N166), .B0(N627), .C0(N708), .Y(N829) );
  OAI22X1TF U826 ( .A0(N221), .A1(N685), .B0(N684), .B1(N277), .Y(N686) );
  AOI21X1TF U827 ( .A0(N302), .A1(N221), .B0(N683), .Y(N684) );
  INVX2TF U828 ( .A(N297), .Y(N821) );
  AOI221X1TF U829 ( .A0(N302), .A1(N277), .B0(N421), .B1(REG_A[13]), .C0(N881), 
        .Y(N685) );
  INVX2TF U830 ( .A(N838), .Y(N881) );
  OAI211X1TF U831 ( .A0(N355), .A1(N267), .B0(N354), .C0(N353), .Y(N356) );
  AND2X2TF U832 ( .A(N422), .B(N424), .Y(N421) );
  NOR2X1TF U833 ( .A(N943), .B(N893), .Y(N953) );
  AOI21X1TF U834 ( .A0(N426), .A1(N422), .B0(N432), .Y(N591) );
  INVX2TF U835 ( .A(N423), .Y(N970) );
  NOR2X2TF U836 ( .A(N304), .B(N169), .Y(N422) );
  AOI31X1TF U837 ( .A0(N854), .A1(N407), .A2(N869), .B0(N351), .Y(N354) );
  AOI22X1TF U838 ( .A0(N706), .A1(N406), .B0(N297), .B1(N349), .Y(N350) );
  OAI21X1TF U839 ( .A0(N843), .A1(N277), .B0(N348), .Y(N349) );
  AOI21X1TF U840 ( .A0(N676), .A1(REG_A[14]), .B0(N623), .Y(N348) );
  NOR2X1TF U841 ( .A(N166), .B(N276), .Y(N623) );
  AND2X2TF U842 ( .A(N407), .B(N428), .Y(N406) );
  INVX2TF U843 ( .A(N595), .Y(N428) );
  AND2X2TF U844 ( .A(N407), .B(N867), .Y(N404) );
  NOR2X2TF U845 ( .A(N211), .B(REG_B[2]), .Y(N867) );
  OAI211X1TF U846 ( .A0(N1014), .A1(N166), .B0(N588), .C0(N692), .Y(N854) );
  INVX2TF U847 ( .A(N842), .Y(N676) );
  AOI21X1TF U848 ( .A0(N420), .A1(N223), .B0(N369), .Y(N355) );
  INVX2TF U849 ( .A(N674), .Y(N876) );
  INVX2TF U850 ( .A(N675), .Y(N347) );
  AND2X2TF U851 ( .A(N407), .B(N309), .Y(N405) );
  NOR2X1TF U852 ( .A(REG_B[2]), .B(REG_B[3]), .Y(N309) );
  AND2X2TF U853 ( .A(N380), .B(N426), .Y(N407) );
  INVX2TF U854 ( .A(N879), .Y(N420) );
  OR2X2TF U855 ( .A(N894), .B(N937), .Y(N879) );
  INVX2TF U856 ( .A(N424), .Y(N937) );
  NOR2X1TF U857 ( .A(N416), .B(N312), .Y(N313) );
  OAI21X1TF U858 ( .A0(N584), .A1(N429), .B0(CODE_TYPE[4]), .Y(N311) );
  NOR2X1TF U859 ( .A(N53), .B(N289), .Y(N584) );
  NOR2X1TF U860 ( .A(CODE_TYPE[3]), .B(N310), .Y(N314) );
  OAI21X1TF U861 ( .A0(N161), .A1(N53), .B0(CODE_TYPE[2]), .Y(N582) );
  OAI21X1TF U862 ( .A0(N380), .A1(N934), .B0(N424), .Y(N306) );
  AND2X2TF U863 ( .A(N263), .B(CODE_TYPE[3]), .Y(N424) );
  AND2X2TF U864 ( .A(N693), .B(N429), .Y(N380) );
  INVX2TF U865 ( .A(N940), .Y(N305) );
  OAI22X1TF U866 ( .A0(N800), .A1(N172), .B0(N300), .B1(N59), .Y(N1007) );
  OAI22X1TF U867 ( .A0(N799), .A1(N172), .B0(N300), .B1(N271), .Y(N1001) );
  OAI22X1TF U868 ( .A0(N794), .A1(N172), .B0(N300), .B1(N272), .Y(N957) );
  OAI22X1TF U869 ( .A0(N798), .A1(N172), .B0(N300), .B1(N273), .Y(N994) );
  OAI22X1TF U870 ( .A0(N796), .A1(N172), .B0(N300), .B1(N282), .Y(N979) );
  OAI22X1TF U871 ( .A0(N787), .A1(N172), .B0(N300), .B1(N278), .Y(N1212) );
  OAI22X1TF U872 ( .A0(N791), .A1(N172), .B0(N300), .B1(N283), .Y(N1024) );
  OAI22X1TF U873 ( .A0(N793), .A1(N173), .B0(N300), .B1(N274), .Y(N1154) );
  OAI22X1TF U874 ( .A0(N789), .A1(N173), .B0(N300), .B1(N276), .Y(N1188) );
  OAI22X1TF U875 ( .A0(N790), .A1(N173), .B0(N160), .B1(N287), .Y(N1021) );
  OAI22X1TF U876 ( .A0(N788), .A1(N173), .B0(N160), .B1(N277), .Y(N1200) );
  OAI22X1TF U877 ( .A0(N792), .A1(N173), .B0(N160), .B1(N266), .Y(N1173) );
  OAI22X1TF U878 ( .A0(N786), .A1(N173), .B0(N160), .B1(N267), .Y(N1018) );
  OAI22X1TF U879 ( .A0(N797), .A1(N172), .B0(N300), .B1(N280), .Y(N1167) );
  OAI22X1TF U880 ( .A0(N795), .A1(N173), .B0(N160), .B1(N279), .Y(N1160) );
  AOI22X1TF U881 ( .A0(N184), .A1(REG_A[13]), .B0(N862), .B1(REG_A[11]), .Y(
        N705) );
  AOI22X1TF U882 ( .A0(N184), .A1(REG_A[12]), .B0(N862), .B1(REG_A[14]), .Y(
        N866) );
  INVX2TF U883 ( .A(N426), .Y(N969) );
  AOI21X1TF U884 ( .A0(N862), .A1(REG_A[2]), .B0(N611), .Y(N822) );
  AOI22X1TF U885 ( .A0(N184), .A1(REG_A[2]), .B0(N862), .B1(REG_A[4]), .Y(N599) );
  AOI21X1TF U886 ( .A0(N347), .A1(REG_A[13]), .B0(N624), .Y(N688) );
  AOI22X1TF U887 ( .A0(N184), .A1(REG_A[3]), .B0(N862), .B1(REG_A[5]), .Y(N627) );
  NAND2X1TF U888 ( .A(N161), .B(CODE_TYPE[2]), .Y(N304) );
  AOI22X1TF U889 ( .A0(N184), .A1(REG_A[1]), .B0(N862), .B1(REG_A[3]), .Y(N588) );
  AOI21X1TF U890 ( .A0(N347), .A1(N162), .B0(N876), .Y(N715) );
  INVX2TF U891 ( .A(N963), .Y(N492) );
  MXI2X1TF U892 ( .A(N294), .B(N393), .S0(N409), .Y(N448) );
  NAND2X1TF U893 ( .A(N1237), .B(N395), .Y(N391) );
  NAND2X1TF U894 ( .A(N393), .B(N379), .Y(N888) );
  NAND4BX1TF U895 ( .AN(N1175), .B(N400), .C(N401), .D(N377), .Y(N378) );
  OAI2BB1X1TF U896 ( .A0N(N474), .A1N(N159), .B0(N344), .Y(N345) );
  AO21X1TF U897 ( .A0(N159), .A1(N468), .B0(N319), .Y(N698) );
  NAND2X1TF U898 ( .A(N874), .B(N502), .Y(N318) );
  NAND4BX1TF U899 ( .AN(N1184), .B(N402), .C(N409), .D(N399), .Y(N376) );
  NOR2BX1TF U900 ( .AN(N736), .B(N328), .Y(N329) );
  OAI2BB1X1TF U901 ( .A0N(N297), .A1N(N854), .B0(N327), .Y(N328) );
  AO22X1TF U902 ( .A0(N504), .A1(N874), .B0(N709), .B1(N162), .Y(N326) );
  AOI2BB1X1TF U903 ( .A0N(N822), .A1N(N821), .B0(N333), .Y(N334) );
  AO21X1TF U904 ( .A0(N851), .A1(N819), .B0(N332), .Y(N333) );
  OAI2BB1X1TF U905 ( .A0N(N469), .A1N(N159), .B0(N331), .Y(N332) );
  OA21XLTF U906 ( .A0(N828), .A1(N827), .B0(N330), .Y(N331) );
  NAND2X1TF U907 ( .A(N503), .B(N874), .Y(N330) );
  NAND2BX1TF U908 ( .AN(N836), .B(N342), .Y(N1175) );
  NAND3X1TF U909 ( .A(N340), .B(N339), .C(N338), .Y(N341) );
  NAND2X1TF U910 ( .A(N337), .B(REG_B[9]), .Y(N340) );
  NAND2X1TF U911 ( .A(N204), .B(N336), .Y(N337) );
  AOI2BB2X1TF U912 ( .B0(N295), .B1(REG_A[9]), .A0N(N879), .A1N(REG_A[9]), .Y(
        N336) );
  NAND2X1TF U913 ( .A(N398), .B(IO_DATAINB[0]), .Y(N386) );
  NAND2X1TF U914 ( .A(N421), .B(REG_A[0]), .Y(N368) );
  NAND2X1TF U915 ( .A(N477), .B(N180), .Y(N365) );
  AOI2BB2X1TF U916 ( .B0(N668), .B1(N297), .A0N(N220), .A1N(N672), .Y(N358) );
  NAND2X1TF U917 ( .A(N479), .B(N180), .Y(N362) );
  NAND2BX1TF U918 ( .AN(N687), .B(N323), .Y(N324) );
  CLKBUFX2TF U919 ( .A(N420), .Y(N302) );
  AO21X1TF U920 ( .A0(N204), .A1(N352), .B0(N223), .Y(N353) );
  MXI2X1TF U921 ( .A(N420), .B(N421), .S0(REG_A[15]), .Y(N352) );
  OAI2BB1X1TF U922 ( .A0N(N860), .A1N(N404), .B0(N350), .Y(N351) );
  OAI2BB1X1TF U923 ( .A0N(N297), .A1N(N862), .B0(N715), .Y(N369) );
  CLKBUFX2TF U924 ( .A(N421), .Y(N295) );
  CLKBUFX2TF U925 ( .A(N405), .Y(N297) );
  CLKBUFX2TF U926 ( .A(N420), .Y(N303) );
  NAND3X1TF U927 ( .A(I_ADDR[1]), .B(I_ADDR[2]), .C(I_ADDR[3]), .Y(N566) );
  NAND2X1TF U928 ( .A(N563), .B(I_ADDR[4]), .Y(N562) );
  NOR2BX1TF U929 ( .AN(I_ADDR[5]), .B(N562), .Y(N558) );
  NAND2X1TF U930 ( .A(N558), .B(I_ADDR[6]), .Y(N557) );
  NOR2BX1TF U931 ( .AN(I_ADDR[7]), .B(N557), .Y(N570) );
  NOR2BX1TF U932 ( .AN(N525), .B(N555), .Y(N165) );
  NAND4X1TF U933 ( .A(STATE[2]), .B(N270), .C(N262), .D(N291), .Y(N544) );
  OAI221XLTF U934 ( .A0(N693), .A1(N263), .B0(N289), .B1(N423), .C0(N169), .Y(
        N437) );
  NAND2BX1TF U935 ( .AN(N551), .B(START), .Y(N533) );
  AND4X1TF U936 ( .A(N794), .B(N797), .C(N796), .D(N795), .Y(N539) );
  OAI2BB2XLTF U937 ( .B0(N540), .B1(N535), .A0N(N525), .A1N(N555), .Y(N527) );
  NAND2X1TF U939 ( .A(N263), .B(N429), .Y(N936) );
  NAND2X1TF U940 ( .A(CODE_TYPE[4]), .B(N580), .Y(N941) );
  NAND2X1TF U941 ( .A(N299), .B(REG_A[6]), .Y(N630) );
  NAND2X1TF U942 ( .A(N56), .B(REG_A[4]), .Y(N690) );
  NAND2X1TF U943 ( .A(N183), .B(REG_A[5]), .Y(N707) );
  NAND2X1TF U944 ( .A(REG_A[7]), .B(N862), .Y(N711) );
  NAND4X1TF U945 ( .A(N630), .B(N690), .C(N707), .D(N711), .Y(N860) );
  NAND2X1TF U946 ( .A(REG_A[10]), .B(N299), .Y(N619) );
  NAND2X1TF U947 ( .A(N56), .B(REG_A[8]), .Y(N631) );
  NAND2X1TF U948 ( .A(N184), .B(REG_A[9]), .Y(N710) );
  NAND2X1TF U949 ( .A(N862), .B(REG_A[11]), .Y(N5860) );
  NAND4X1TF U950 ( .A(N619), .B(N631), .C(N710), .D(N5860), .Y(N706) );
  NAND2X1TF U951 ( .A(N211), .B(REG_B[2]), .Y(N595) );
  NAND2X1TF U952 ( .A(N299), .B(REG_A[2]), .Y(N692) );
  NAND3X1TF U953 ( .A(N57), .B(N211), .C(N408), .Y(N827) );
  NAND2X1TF U954 ( .A(N183), .B(REG_A[6]), .Y(N603) );
  NAND2X1TF U955 ( .A(REG_A[8]), .B(N347), .Y(N600) );
  NAND2X1TF U956 ( .A(REG_A[7]), .B(N299), .Y(N612) );
  NAND4BX1TF U957 ( .AN(N737), .B(N603), .C(N600), .D(N612), .Y(N669) );
  NAND2X1TF U958 ( .A(N299), .B(REG_A[13]), .Y(N865) );
  NAND2X1TF U959 ( .A(REG_A[10]), .B(N183), .Y(N666) );
  NAND2X1TF U960 ( .A(N56), .B(REG_A[11]), .Y(N864) );
  NAND4BX1TF U961 ( .AN(N644), .B(N600), .C(N666), .D(N864), .Y(N841) );
  NAND2X1TF U962 ( .A(N299), .B(REG_A[5]), .Y(N607) );
  NAND2X1TF U963 ( .A(N347), .B(REG_A[4]), .Y(N604) );
  NAND4BX1TF U964 ( .AN(N647), .B(N607), .C(N604), .D(N603), .Y(N840) );
  NAND2X1TF U965 ( .A(N867), .B(N408), .Y(N856) );
  NAND2X1TF U966 ( .A(N184), .B(REG_A[4]), .Y(N608) );
  NAND2X1TF U967 ( .A(N347), .B(REG_A[6]), .Y(N615) );
  NAND4BX1TF U968 ( .AN(N845), .B(N608), .C(N607), .D(N615), .Y(N868) );
  NAND2X1TF U969 ( .A(N299), .B(REG_A[11]), .Y(N667) );
  NAND2X1TF U970 ( .A(REG_A[9]), .B(N347), .Y(N677) );
  NAND2X1TF U971 ( .A(N184), .B(REG_A[11]), .Y(N620) );
  NAND4BX1TF U972 ( .AN(N623), .B(N677), .C(N620), .D(N619), .Y(N832) );
  NAND2X1TF U973 ( .A(N299), .B(REG_A[4]), .Y(N708) );
  NAND2X1TF U974 ( .A(N407), .B(N211), .Y(N628) );
  OAI2BB1X1TF U975 ( .A0N(N303), .A1N(N213), .B0(N674), .Y(N635) );
  NAND2X1TF U976 ( .A(REG_A[7]), .B(N183), .Y(N678) );
  NAND2X1TF U977 ( .A(N862), .B(REG_A[5]), .Y(N632) );
  NAND4X1TF U978 ( .A(N678), .B(N632), .C(N631), .D(N630), .Y(N689) );
  NAND4X1TF U979 ( .A(N1178), .B(N1171), .C(N1165), .D(N1162), .Y(N889) );
  AOI2BB2X1TF U980 ( .B0(REG_B[2]), .B1(N652), .A0N(N650), .A1N(REG_B[2]), .Y(
        N653) );
  NAND2X1TF U981 ( .A(N408), .B(N653), .Y(N820) );
  AOI222XLTF U982 ( .A0(N671), .A1(N867), .B0(N869), .B1(N670), .C0(N669), 
        .C1(N428), .Y(N673) );
  NAND2X1TF U983 ( .A(N299), .B(REG_A[12]), .Y(N704) );
  NAND2X1TF U984 ( .A(REG_A[10]), .B(N56), .Y(N712) );
  NAND2X1TF U985 ( .A(N56), .B(REG_A[6]), .Y(N680) );
  NAND2X1TF U986 ( .A(REG_A[8]), .B(N299), .Y(N713) );
  NAND4X1TF U987 ( .A(N680), .B(N678), .C(N713), .D(N677), .Y(N837) );
  NAND2X1TF U988 ( .A(REG_B[3]), .B(N407), .Y(N681) );
  OAI221XLTF U989 ( .A0(REG_A[1]), .A1(N879), .B0(N59), .B1(N880), .C0(N838), 
        .Y(N700) );
  NAND2X1TF U990 ( .A(N694), .B(N57), .Y(N834) );
  NAND4X1TF U991 ( .A(N713), .B(N712), .C(N711), .D(N710), .Y(N853) );
  AOI2BB2X1TF U992 ( .B0(REG_A[3]), .B1(N718), .A0N(N211), .A1N(N717), .Y(N719) );
  OAI2BB2XLTF U993 ( .B0(N830), .B1(N266), .A0N(N510), .A1N(N874), .Y(N836) );
  OAI2BB2XLTF U994 ( .B0(N852), .B1(N272), .A0N(N508), .A1N(N874), .Y(N859) );
  NAND2X1TF U995 ( .A(N57), .B(N211), .Y(N863) );
  AO22X1TF U996 ( .A0(N870), .A1(N869), .B0(N868), .B1(N867), .Y(N871) );
  AOI2BB1X1TF U997 ( .A0N(N429), .A1N(N934), .B0(N969), .Y(N895) );
  NAND2X1TF U998 ( .A(CODE_TYPE[3]), .B(N940), .Y(N892) );
  NAND2X1TF U999 ( .A(N961), .B(N917), .Y(N974) );
  NAND2X1TF U1000 ( .A(N426), .B(N934), .Y(N935) );
  NOR2X1TF U1001 ( .A(N950), .B(N281), .Y(N945) );
  NAND2X1TF U1002 ( .A(N947), .B(N412), .Y(N946) );
  NAND2X1TF U1003 ( .A(N947), .B(N281), .Y(N949) );
  NAND2X1TF U1004 ( .A(N260), .B(N275), .Y(N962) );
  AOI2BB2X1TF U1005 ( .B0(IO_DATAINA[5]), .B1(N298), .A0N(N1162), .A1N(N1225), 
        .Y(N972) );
  AOI2BB2X1TF U1006 ( .B0(IO_DATAINB[10]), .B1(N398), .A0N(N410), .A1N(N427), 
        .Y(N1139) );
  AOI2BB2X1TF U1007 ( .B0(IO_DATAINB[8]), .B1(N398), .A0N(N410), .A1N(N425), 
        .Y(N1158) );
  AOI2BB2X1TF U1008 ( .B0(IO_DATAINA[6]), .B1(N298), .A0N(N1162), .A1N(N1224), 
        .Y(N1163) );
  AOI2BB2X1TF U1009 ( .B0(IO_DATAINB[9]), .B1(N398), .A0N(N410), .A1N(N419), 
        .Y(N1177) );
  AOI2BB2X1TF U1010 ( .B0(IO_DATAINB[12]), .B1(N398), .A0N(N410), .A1N(N418), 
        .Y(N1191) );
  AOI2BB2X1TF U1011 ( .B0(IO_DATAINB[11]), .B1(N398), .A0N(N410), .A1N(N415), 
        .Y(N1198) );
  OAI2BB1X1TF U1012 ( .A0N(N1223), .A1N(N396), .B0(N1203), .Y(N629) );
  NAND2X1TF U1013 ( .A(N1217), .B(N1216), .Y(N637) );
endmodule


module SCPU_SRAM_8BIT_ALU_SPI_TOP_VG ( CLK, RST_N, CTRL_MODE, CTRL_BGN, CPU_BGN, 
        LOAD_N, CTRL_SI, ADC_PI, CTRL_RDY, CTRL_SO, NXT, SCLK1, SCLK2, LAT, 
        SPI_SO );
  input [1:0] CTRL_MODE;
  input [15:0] ADC_PI;
  output [1:0] NXT;
  input CLK, RST_N, CTRL_BGN, CPU_BGN, LOAD_N, CTRL_SI;
  output CTRL_RDY, CTRL_SO, SCLK1, SCLK2, LAT, SPI_SO;
  wire   CEN_AFTER_MUX, WEN_AFTER_MUX, I_CLK, I_RST_N, I_CTRL_BGN, I_CPU_BGN,
         I_LOAD_N, I_CTRL_SI, I_CTRL_SO, I_SCLK1, I_SCLK2, I_SPI_SO,
         SCPU_CTRL_SPI_CEN, \SCPU_CTRL_SPI_IO_DATAOUTB[0] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[1] , \SCPU_CTRL_SPI_IO_DATAOUTB[2] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[3] , \SCPU_CTRL_SPI_IO_DATAOUTB[4] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[5] , \SCPU_CTRL_SPI_IO_DATAOUTB[6] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[7] , \SCPU_CTRL_SPI_IO_DATAOUTB[8] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[9] , \SCPU_CTRL_SPI_IO_DATAOUTB[10] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[11] , \SCPU_CTRL_SPI_IO_DATAOUTB[12] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[0] , \SCPU_CTRL_SPI_IO_DATAOUTA[1] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[2] , \SCPU_CTRL_SPI_IO_DATAOUTA[3] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[4] , \SCPU_CTRL_SPI_IO_DATAOUTA[5] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[6] , \SCPU_CTRL_SPI_IO_DATAOUTA[7] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[8] , \SCPU_CTRL_SPI_IO_DATAOUTA[9] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[10] , \SCPU_CTRL_SPI_IO_DATAOUTA[11] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[12] , \SCPU_CTRL_SPI_IO_CONTROL[0] ,
         \SCPU_CTRL_SPI_IO_CONTROL[1] , \SCPU_CTRL_SPI_IO_CONTROL[2] ,
         \SCPU_CTRL_SPI_IO_CONTROL[3] , \SCPU_CTRL_SPI_IO_CONTROL[4] ,
         \SCPU_CTRL_SPI_IO_CONTROL[5] , \SCPU_CTRL_SPI_IO_CONTROL[6] ,
         SCPU_CTRL_SPI_D_WE, SCPU_CTRL_SPI_IS_I_ADDR, SCPU_CTRL_SPI_CCT_N54,
         SCPU_CTRL_SPI_CCT_N53, SCPU_CTRL_SPI_CCT_N51, SCPU_CTRL_SPI_CCT_N50,
         SCPU_CTRL_SPI_CCT_N49, SCPU_CTRL_SPI_CCT_N24,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] , \SCPU_CTRL_SPI_CCT_REG_BITS[1] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[2] , \SCPU_CTRL_SPI_CCT_REG_BITS[3] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[4] , \SCPU_CTRL_SPI_CCT_REG_BITS[5] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[6] , \SCPU_CTRL_SPI_CCT_REG_BITS[7] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[8] , \SCPU_CTRL_SPI_CCT_REG_BITS[9] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[10] , \SCPU_CTRL_SPI_CCT_REG_BITS[11] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[12] , \SCPU_CTRL_SPI_CCT_REG_BITS[13] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[14] , \SCPU_CTRL_SPI_CCT_REG_BITS[15] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[16] , \SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ,
         SCPU_CTRL_SPI_PUT_N108, SCPU_CTRL_SPI_PUT_N107,
         SCPU_CTRL_SPI_PUT_N106, \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ,
         \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ,
         \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ,
         \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] , \SCPU_CTRL_SPI_PUT_SPI_STATE[0] ,
         \SCPU_CTRL_SPI_PUT_SPI_STATE[1] , \SCPU_CTRL_SPI_PUT_CNT_STATE[1] ,
         \SCPU_CTRL_SPI_PUT_CNT_STATE[2] , N31, N32, N33, N34, N35, N36, N37,
         N38, N39, N40, N41, N42, N43, N44, N45, N78, N79, N80, N81, N82, N83,
         N84, N85, N86, N91, N93, N100, N102, N103, N158, N189, N190, N191,
         N192, N193, N194, N195, N196, N197, N198, N199, N200, N201, N202,
         N203, N204, N205, N206, N207, N208, N209, N210, N212, N213, N214,
         N215, N216, N218, N219, N220, N221, N222, N233, N234, N241, N267,
         N268, N269, N270, N271, N272, N273, N278, N279, N280, N281, N282,
         N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293,
         N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304,
         N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315,
         N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326,
         N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337,
         N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, N348,
         N349, N350, N351, N352, N353, N354, N355, N356, N357, N358, N359,
         N360, N361, N362, N363, N364, N365, N366, N367, N368, N369, N370,
         N371, N372, N373, N374, N375, N376, N377, N378, N379, N380, N381,
         N382, N383, N384, N385, N386, N387, N388, N389, N390, N391, N392,
         N393, N394, N395, N396, N397, N398, N399, N400, N401, N402, N403,
         N404, N405, N406, N407, N408, N409, N410, N411, N412, N413, N414,
         N415, N416, N417, N418, N419, N420, N421, N422, N423, N424, N425,
         N426, N427, N428, N429;
  wire   [8:0] A_AFTER_MUX;
  wire   [7:0] D_AFTER_MUX;
  wire   [7:0] Q_FROM_SRAM;
  wire   [1:0] I_CTRL_MODE;
  wire   [15:0] I_ADC_PI;
  wire   [1:0] I_NXT;
  wire   [8:0] SCPU_CTRL_SPI_A_SPI;
  wire   [12:0] SCPU_CTRL_SPI_POUT;
  wire   [12:0] SCPU_CTRL_SPI_FOUT;
  wire   [9:0] SCPU_CTRL_SPI_IO_OFFSET;
  wire   [15:0] SCPU_CTRL_SPI_IO_DATAINA;
  wire   [0:0] SCPU_CTRL_SPI_IO_STATUS;
  wire   [7:0] SCPU_CTRL_SPI_D_DATAOUT;
  wire   [8:1] SCPU_CTRL_SPI_D_ADDR;
  wire   [8:0] SCPU_CTRL_SPI_I_ADDR;
  wire   [7:0] SCPU_CTRL_SPI_D_DATAIN;
  wire   [7:0] SCPU_CTRL_SPI_I_DATAIN;
  wire   [7:1] SCPU_CTRL_SPI_PUT_SRAM_REGS;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21;

  RA1SHD_IBM512X8 sram ( .Q(Q_FROM_SRAM), .A(A_AFTER_MUX), .D(D_AFTER_MUX), 
        .CLK(I_CLK), .CEN(CEN_AFTER_MUX), .WEN(WEN_AFTER_MUX) );
  PIC ipad_clk ( .IE(1'b1), .P(CLK), .Y(I_CLK) );
  PIC ipad_rst_n ( .IE(1'b1), .P(RST_N), .Y(I_RST_N) );
  PIC ipad_ctrl_mode0 ( .IE(1'b1), .P(CTRL_MODE[0]), .Y(I_CTRL_MODE[0]) );
  PIC ipad_ctrl_mode1 ( .IE(1'b1), .P(CTRL_MODE[1]), .Y(I_CTRL_MODE[1]) );
  PIC ipad_ctrl_bgn ( .IE(1'b1), .P(CTRL_BGN), .Y(I_CTRL_BGN) );
  PIC ipad_cpu_str ( .IE(1'b1), .P(CPU_BGN), .Y(I_CPU_BGN) );
  PIC ipad_load_n ( .IE(1'b1), .P(LOAD_N), .Y(I_LOAD_N) );
  PIC ipad_ctrl_si ( .IE(1'b1), .P(CTRL_SI), .Y(I_CTRL_SI) );
  PIC ipad_adc_pi0 ( .IE(1'b1), .P(ADC_PI[0]), .Y(I_ADC_PI[0]) );
  PIC ipad_adc_pi1 ( .IE(1'b1), .P(ADC_PI[1]), .Y(I_ADC_PI[1]) );
  PIC ipad_adc_pi2 ( .IE(1'b1), .P(ADC_PI[2]), .Y(I_ADC_PI[2]) );
  PIC ipad_adc_pi3 ( .IE(1'b1), .P(ADC_PI[3]), .Y(I_ADC_PI[3]) );
  PIC ipad_adc_pi4 ( .IE(1'b1), .P(ADC_PI[4]), .Y(I_ADC_PI[4]) );
  PIC ipad_adc_pi5 ( .IE(1'b1), .P(ADC_PI[5]), .Y(I_ADC_PI[5]) );
  PIC ipad_adc_pi6 ( .IE(1'b1), .P(ADC_PI[6]), .Y(I_ADC_PI[6]) );
  PIC ipad_adc_pi7 ( .IE(1'b1), .P(ADC_PI[7]), .Y(I_ADC_PI[7]) );
  PIC ipad_adc_pi8 ( .IE(1'b1), .P(ADC_PI[8]), .Y(I_ADC_PI[8]) );
  PIC ipad_adc_pi9 ( .IE(1'b1), .P(ADC_PI[9]), .Y(I_ADC_PI[9]) );
  PIC ipad_adc_pi10 ( .IE(1'b1), .P(ADC_PI[10]), .Y(I_ADC_PI[10]) );
  PIC ipad_adc_pi11 ( .IE(1'b1), .P(ADC_PI[11]), .Y(I_ADC_PI[11]) );
  PIC ipad_adc_pi12 ( .IE(1'b1), .P(ADC_PI[12]), .Y(I_ADC_PI[12]) );
  PIC ipad_adc_pi13 ( .IE(1'b1), .P(ADC_PI[13]), .Y(I_ADC_PI[13]) );
  PIC ipad_adc_pi14 ( .IE(1'b1), .P(ADC_PI[14]), .Y(I_ADC_PI[14]) );
  PIC ipad_adc_pi15 ( .IE(1'b1), .P(ADC_PI[15]), .Y(I_ADC_PI[15]) );
  POC8B opad_ctrl_rdy ( .A(N220), .P(CTRL_RDY) );
  POC8B opad_ctrl_so ( .A(I_CTRL_SO), .P(CTRL_SO) );
  POC8B opad_nxt0 ( .A(I_NXT[0]), .P(NXT[0]) );
  POC8B opad_nxt1 ( .A(I_NXT[1]), .P(NXT[1]) );
  POC8B opad_sclk1 ( .A(I_SCLK1), .P(SCLK1) );
  POC8B opad_sclk2 ( .A(I_SCLK2), .P(SCLK2) );
  POC8B opad_lat ( .A(N222), .P(LAT) );
  POC8B opad_spi_so ( .A(I_SPI_SO), .P(SPI_SO) );
  SHARE_SUPERALU_VG \scpu_ctrl_spi/ALU_01  ( .CLK(I_CLK), .RST_N(I_RST_N), .X_IN(
        {\SCPU_CTRL_SPI_IO_DATAOUTA[12] , \SCPU_CTRL_SPI_IO_DATAOUTA[11] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[10] , \SCPU_CTRL_SPI_IO_DATAOUTA[9] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[8] , \SCPU_CTRL_SPI_IO_DATAOUTA[7] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[6] , \SCPU_CTRL_SPI_IO_DATAOUTA[5] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[4] , \SCPU_CTRL_SPI_IO_DATAOUTA[3] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[2] , \SCPU_CTRL_SPI_IO_DATAOUTA[1] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[0] }), .Y_IN({
        \SCPU_CTRL_SPI_IO_DATAOUTB[12] , \SCPU_CTRL_SPI_IO_DATAOUTB[11] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[10] , \SCPU_CTRL_SPI_IO_DATAOUTB[9] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[8] , \SCPU_CTRL_SPI_IO_DATAOUTB[7] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[6] , \SCPU_CTRL_SPI_IO_DATAOUTB[5] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[4] , \SCPU_CTRL_SPI_IO_DATAOUTB[3] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[2] , \SCPU_CTRL_SPI_IO_DATAOUTB[1] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[0] }), .ALU_START(
        \SCPU_CTRL_SPI_IO_CONTROL[5] ), .ALU_TYPE({
        \SCPU_CTRL_SPI_IO_CONTROL[4] , \SCPU_CTRL_SPI_IO_CONTROL[3] , 
        \SCPU_CTRL_SPI_IO_CONTROL[2] }), .MODE_TYPE({
        \SCPU_CTRL_SPI_IO_CONTROL[1] , \SCPU_CTRL_SPI_IO_CONTROL[0] }), 
        .OFFSET(SCPU_CTRL_SPI_IO_OFFSET), .FOUT(SCPU_CTRL_SPI_FOUT), .POUT(
        SCPU_CTRL_SPI_POUT), .ALU_IS_DONE(SCPU_CTRL_SPI_IO_STATUS[0]) );
  SERIAL_CPU_8BIT_VG \scpu_ctrl_spi/uut  ( .CLK(I_CLK), .ENABLE(1'b0), .RST_N(
        I_RST_N), .START(I_CPU_BGN), .I_DATAIN(SCPU_CTRL_SPI_I_DATAIN), 
        .D_DATAIN(SCPU_CTRL_SPI_D_DATAIN), .IS_I_ADDR(SCPU_CTRL_SPI_IS_I_ADDR), 
        .NXT(I_NXT), .I_ADDR(SCPU_CTRL_SPI_I_ADDR), .D_ADDR({
        SCPU_CTRL_SPI_D_ADDR, SYNOPSYS_UNCONNECTED__0}), .D_WE(
        SCPU_CTRL_SPI_D_WE), .D_DATAOUT(SCPU_CTRL_SPI_D_DATAOUT), .IO_STATUS({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, N221, SCPU_CTRL_SPI_IO_STATUS[0]}), .IO_CONTROL({
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, \SCPU_CTRL_SPI_IO_CONTROL[6] , 
        \SCPU_CTRL_SPI_IO_CONTROL[5] , \SCPU_CTRL_SPI_IO_CONTROL[4] , 
        \SCPU_CTRL_SPI_IO_CONTROL[3] , \SCPU_CTRL_SPI_IO_CONTROL[2] , 
        \SCPU_CTRL_SPI_IO_CONTROL[1] , \SCPU_CTRL_SPI_IO_CONTROL[0] }), 
        .IO_DATAINA(SCPU_CTRL_SPI_IO_DATAINA), .IO_DATAINB({1'b0, 1'b0, 1'b0, 
        SCPU_CTRL_SPI_POUT}), .IO_DATAOUTA({SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        \SCPU_CTRL_SPI_IO_DATAOUTA[12] , \SCPU_CTRL_SPI_IO_DATAOUTA[11] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[10] , \SCPU_CTRL_SPI_IO_DATAOUTA[9] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[8] , \SCPU_CTRL_SPI_IO_DATAOUTA[7] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[6] , \SCPU_CTRL_SPI_IO_DATAOUTA[5] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[4] , \SCPU_CTRL_SPI_IO_DATAOUTA[3] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[2] , \SCPU_CTRL_SPI_IO_DATAOUTA[1] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[0] }), .IO_DATAOUTB({
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, \SCPU_CTRL_SPI_IO_DATAOUTB[12] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[11] , \SCPU_CTRL_SPI_IO_DATAOUTB[10] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[9] , \SCPU_CTRL_SPI_IO_DATAOUTB[8] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[7] , \SCPU_CTRL_SPI_IO_DATAOUTB[6] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[5] , \SCPU_CTRL_SPI_IO_DATAOUTB[4] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[3] , \SCPU_CTRL_SPI_IO_DATAOUTB[2] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[1] , \SCPU_CTRL_SPI_IO_DATAOUTB[0] }), 
        .IO_OFFSET({SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SCPU_CTRL_SPI_IO_OFFSET}) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[5]  ( .D(N158), .RN(
        SCPU_CTRL_SPI_CCT_N53), .CK(I_CLK), .QN(N288) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[3]  ( .D(N158), .RN(
        SCPU_CTRL_SPI_CCT_N51), .CK(I_CLK), .QN(N287) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[2]  ( .D(N158), .RN(
        SCPU_CTRL_SPI_CCT_N50), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[1]  ( .D(N158), .RN(
        SCPU_CTRL_SPI_CCT_N49), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[6]  ( .D(N158), .RN(
        SCPU_CTRL_SPI_CCT_N54), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[4]  ( .D(N45), .CK(I_CLK), 
        .SN(N44), .RN(N43), .QN(N284) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[0]  ( .D(N33), .CK(I_CLK), 
        .SN(N32), .RN(N31), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .QN(N283)
         );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[3]  ( .D(N42), .CK(I_CLK), 
        .SN(N41), .RN(N40), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] ), .QN(N281)
         );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[2]  ( .D(N39), .CK(I_CLK), 
        .SN(N38), .RN(N37), .QN(N280) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[1]  ( .D(N36), .CK(I_CLK), 
        .SN(N35), .RN(N34), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ), .QN(N278)
         );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[7]  ( .D(N204), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[7]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[6]  ( .D(N198), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[6]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[5]  ( .D(N199), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[5]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[4]  ( .D(N200), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[4]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[3]  ( .D(N201), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[3]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[2]  ( .D(N202), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[2]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[1]  ( .D(N203), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[1]) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[7]  ( .D(N189), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[7] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[6]  ( .D(N190), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[6] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[5]  ( .D(N191), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[5] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[4]  ( .D(N192), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[4] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[3]  ( .D(N193), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[3] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[2]  ( .D(N194), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[2] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[1]  ( .D(N195), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[1] ) );
  DFFRX2TF \scpu_ctrl_spi/put/cnt_state_reg[2]  ( .D(SCPU_CTRL_SPI_PUT_N108), 
        .CK(I_CLK), .RN(N267), .Q(\SCPU_CTRL_SPI_PUT_CNT_STATE[2] ) );
  DFFRX2TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[2]  ( .D(N207), .CK(I_CLK), 
        .RN(N267), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ) );
  DFFRX2TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[1]  ( .D(N206), .CK(I_CLK), 
        .RN(N267), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[0]  ( .D(N197), .CK(I_CLK), .Q(
        I_SPI_SO) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[0]  ( .D(N196), .CK(I_CLK), .Q(
        I_CTRL_SO) );
  DFFQX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[4]  ( .D(N215), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ) );
  DFFSX2TF \scpu_ctrl_spi/put/cnt_state_reg[0]  ( .D(SCPU_CTRL_SPI_PUT_N106), 
        .CK(I_CLK), .SN(N268), .Q(N290), .QN(N102) );
  DFFQX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[0]  ( .D(N214), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ) );
  DFFRX2TF \scpu_ctrl_spi/put/spi_state_reg[0]  ( .D(N209), .CK(I_CLK), .RN(
        N267), .Q(\SCPU_CTRL_SPI_PUT_SPI_STATE[0] ) );
  DFFRX1TF \scpu_ctrl_spi/put/cnt_state_reg[1]  ( .D(SCPU_CTRL_SPI_PUT_N107), 
        .CK(I_CLK), .RN(N268), .Q(\SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .QN(N286)
         );
  DFFNSRX4TF \scpu_ctrl_spi/put/spi_MUX_reg  ( .D(N213), .CKN(I_CLK), .SN(1'b1), .RN(1'b1), .Q(N279), .QN(N103) );
  DFFNSRXLTF \scpu_ctrl_spi/cct/D_WE_reg  ( .D(N218), .CKN(I_CLK), .SN(1'b1), 
        .RN(1'b1), .QN(N93) );
  DFFNSRX1TF \scpu_ctrl_spi/put/sram_addr_reg[7]  ( .D(N85), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[7]), .QN(N291) );
  DFFNSRXLTF \scpu_ctrl_spi/cct/CEN_reg  ( .D(N219), .CKN(I_CLK), .SN(1'b1), 
        .RN(1'b1), .Q(SCPU_CTRL_SPI_CEN) );
  DFFNSRXLTF \scpu_ctrl_spi/put/sram_addr_reg[8]  ( .D(N86), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[8]) );
  DFFX1TF \scpu_ctrl_spi/cct/ctrl_state_reg[0]  ( .D(N216), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .QN(N368) );
  EDFFTRXLTF \scpu_ctrl_spi/cct/ctrl_state_reg[1]  ( .RN(I_CTRL_BGN), .D(1'b1), 
        .E(N234), .CK(I_CLK), .Q(N285), .QN(N91) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[16]  ( .D(I_CTRL_SI), .E(N241), 
        .CK(I_CLK), .Q(\SCPU_CTRL_SPI_CCT_REG_BITS[16] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[15]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[16] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[15] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[14]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[15] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[14] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[13]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[14] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[13] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[12]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[13] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[12] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[11]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[12] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[11] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[10]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[11] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[10] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[9]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[10] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[9] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[8]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[9] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[8] ) );
  DFFRX2TF \scpu_ctrl_spi/put/spi_state_reg[2]  ( .D(N212), .CK(I_CLK), .RN(
        N268), .Q(N289), .QN(N100) );
  DFFRX2TF \scpu_ctrl_spi/put/spi_state_reg[1]  ( .D(N210), .CK(I_CLK), .RN(
        N267), .Q(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .QN(N282) );
  DFFRX2TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[0]  ( .D(N205), .CK(I_CLK), 
        .RN(N268), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .QN(N292) );
  DFFRX2TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[3]  ( .D(N208), .CK(I_CLK), 
        .RN(N268), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ), .QN(N294) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[1]  ( .D(N79), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[1]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[5]  ( .D(N83), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[5]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[3]  ( .D(N81), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[3]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[2]  ( .D(N80), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[2]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[4]  ( .D(N82), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[4]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[6]  ( .D(N84), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[6]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[0]  ( .D(N78), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[0]), .QN(N293) );
  OR2X2TF U246 ( .A(SCPU_CTRL_SPI_IS_I_ADDR), .B(I_CTRL_BGN), .Y(N381) );
  NOR3X1TF U247 ( .A(N285), .B(\SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .C(N270), 
        .Y(N326) );
  AO21X1TF U248 ( .A0(N278), .A1(N425), .B0(N280), .Y(N233) );
  OAI21X1TF U249 ( .A0(N427), .A1(N428), .B0(N233), .Y(N39) );
  INVX2TF U250 ( .A(N302), .Y(N369) );
  OA21XLTF U251 ( .A0(\SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .A1(I_CTRL_MODE[0]), 
        .B0(N325), .Y(N234) );
  INVX2TF U252 ( .A(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .Y(N295) );
  CLKBUFX2TF U253 ( .A(SCPU_CTRL_SPI_CCT_N24), .Y(N241) );
  AO21XLTF U267 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ), .A1(N299), .B0(
        N300), .Y(SCPU_CTRL_SPI_CCT_N50) );
  OR2X1TF U268 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ), .B(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .Y(N299) );
  OAI21XLTF U269 ( .A0(N380), .A1(N387), .B0(N376), .Y(N191) );
  OAI21XLTF U270 ( .A0(N380), .A1(N388), .B0(N377), .Y(N190) );
  OAI21XLTF U271 ( .A0(N380), .A1(N390), .B0(N379), .Y(N189) );
  OAI21XLTF U272 ( .A0(N380), .A1(N386), .B0(N375), .Y(N192) );
  OAI21XLTF U273 ( .A0(N382), .A1(N380), .B0(N371), .Y(N196) );
  OAI21XLTF U274 ( .A0(N380), .A1(N383), .B0(N372), .Y(N195) );
  OAI21XLTF U275 ( .A0(N380), .A1(N384), .B0(N373), .Y(N194) );
  OAI21XLTF U276 ( .A0(N380), .A1(N385), .B0(N374), .Y(N193) );
  OAI21XLTF U277 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .A1(N332), .B0(
        N331), .Y(N214) );
  NOR3X1TF U278 ( .A(N302), .B(N285), .C(N368), .Y(SCPU_CTRL_SPI_CCT_N24) );
  AOI32X1TF U279 ( .A0(SCPU_CTRL_SPI_A_SPI[0]), .A1(N267), .A2(N427), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[0] ), .B1(N297), .Y(N421) );
  AO21XLTF U280 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ), .A1(N301), .B0(
        N302), .Y(SCPU_CTRL_SPI_CCT_N54) );
  OAI21XLTF U281 ( .A0(N327), .A1(N288), .B0(N301), .Y(SCPU_CTRL_SPI_CCT_N53)
         );
  NAND2XLTF U282 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[4] ), .B(N297), .Y(N44) );
  INVX1TF U283 ( .A(N405), .Y(N408) );
  OAI21XLTF U284 ( .A0(N300), .A1(N287), .B0(N328), .Y(SCPU_CTRL_SPI_CCT_N51)
         );
  NOR2X4TF U285 ( .A(SCPU_CTRL_SPI_CEN), .B(N269), .Y(N323) );
  NAND2XLTF U286 ( .A(N335), .B(N392), .Y(N334) );
  INVX2TF U287 ( .A(I_CTRL_BGN), .Y(N269) );
  NAND2XLTF U288 ( .A(SCPU_CTRL_SPI_A_SPI[0]), .B(SCPU_CTRL_SPI_A_SPI[1]), .Y(
        N418) );
  CLKBUFX2TF U289 ( .A(\SCPU_CTRL_SPI_IO_CONTROL[6] ), .Y(N267) );
  CLKBUFX2TF U290 ( .A(\SCPU_CTRL_SPI_IO_CONTROL[6] ), .Y(N268) );
  INVX2TF U291 ( .A(I_CTRL_BGN), .Y(N270) );
  INVX2TF U292 ( .A(N295), .Y(N271) );
  INVX2TF U293 ( .A(N295), .Y(N272) );
  CLKBUFX2TF U294 ( .A(N241), .Y(N296) );
  NOR3X4TF U295 ( .A(N356), .B(N355), .C(N423), .Y(N365) );
  NOR3X2TF U296 ( .A(\SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .B(
        \SCPU_CTRL_SPI_PUT_CNT_STATE[2] ), .C(N290), .Y(N392) );
  INVX2TF U297 ( .A(N427), .Y(N273) );
  NOR2BX1TF U298 ( .AN(N339), .B(N426), .Y(N424) );
  NAND2X2TF U299 ( .A(SCPU_CTRL_SPI_IS_I_ADDR), .B(N269), .Y(N389) );
  NOR2X1TF U300 ( .A(N390), .B(N381), .Y(SCPU_CTRL_SPI_D_DATAIN[7]) );
  NOR2X1TF U301 ( .A(N388), .B(N381), .Y(SCPU_CTRL_SPI_D_DATAIN[6]) );
  NOR2X1TF U302 ( .A(N386), .B(N381), .Y(SCPU_CTRL_SPI_D_DATAIN[4]) );
  NOR2X1TF U303 ( .A(N384), .B(N381), .Y(SCPU_CTRL_SPI_D_DATAIN[2]) );
  NOR2X1TF U304 ( .A(N383), .B(N381), .Y(SCPU_CTRL_SPI_D_DATAIN[1]) );
  NOR2X1TF U305 ( .A(N387), .B(N381), .Y(SCPU_CTRL_SPI_D_DATAIN[5]) );
  NOR2X1TF U306 ( .A(N385), .B(N381), .Y(SCPU_CTRL_SPI_D_DATAIN[3]) );
  NOR2X1TF U307 ( .A(N382), .B(N381), .Y(SCPU_CTRL_SPI_D_DATAIN[0]) );
  NOR2X1TF U308 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ), .B(N301), .Y(N302)
         );
  NAND2X1TF U309 ( .A(N288), .B(N327), .Y(N301) );
  NOR2X1TF U310 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ), .B(N328), .Y(N327)
         );
  CLKBUFX2TF U311 ( .A(N423), .Y(N297) );
  NOR2X1TF U312 ( .A(N343), .B(N357), .Y(N354) );
  NAND2X1TF U313 ( .A(N369), .B(I_CTRL_BGN), .Y(N332) );
  NAND2X1TF U314 ( .A(N287), .B(N300), .Y(N328) );
  NAND2X1TF U315 ( .A(N333), .B(N100), .Y(N426) );
  NAND2X1TF U316 ( .A(N322), .B(N321), .Y(A_AFTER_MUX[8]) );
  NAND2X1TF U317 ( .A(N317), .B(N316), .Y(A_AFTER_MUX[7]) );
  NAND2X1TF U318 ( .A(N315), .B(N314), .Y(A_AFTER_MUX[6]) );
  NAND2X1TF U319 ( .A(N313), .B(N312), .Y(A_AFTER_MUX[5]) );
  NAND2X1TF U320 ( .A(N311), .B(N310), .Y(A_AFTER_MUX[4]) );
  NAND2X1TF U321 ( .A(N309), .B(N308), .Y(A_AFTER_MUX[3]) );
  NAND2X1TF U322 ( .A(N307), .B(N306), .Y(A_AFTER_MUX[2]) );
  NAND2X1TF U323 ( .A(N305), .B(N304), .Y(A_AFTER_MUX[1]) );
  NOR2X2TF U324 ( .A(N381), .B(N279), .Y(N320) );
  NOR2X2TF U325 ( .A(N279), .B(N389), .Y(N318) );
  NOR2X1TF U326 ( .A(N341), .B(N100), .Y(N355) );
  OR2XLTF U327 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[2] ), .B(N268), .Y(N37) );
  OR2XLTF U328 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[1] ), .B(N268), .Y(N34) );
  OR2XLTF U329 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[3] ), .B(N268), .Y(N40) );
  OR2XLTF U330 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[0] ), .B(N268), .Y(N31) );
  OR2XLTF U331 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[4] ), .B(N268), .Y(N43) );
  OAI2BB2XLTF U332 ( .B0(N395), .B1(N394), .A0N(
        \SCPU_CTRL_SPI_PUT_CNT_STATE[2] ), .A1N(N393), .Y(
        SCPU_CTRL_SPI_PUT_N108) );
  NOR2X1TF U333 ( .A(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ), .B(N338), .Y(N343)
         );
  OAI2BB2XLTF U334 ( .B0(N368), .B1(N332), .A0N(N326), .A1N(N325), .Y(N216) );
  NOR2BX1TF U335 ( .AN(N342), .B(N100), .Y(N222) );
  OAI2BB1X1TF U336 ( .A0N(\SCPU_CTRL_SPI_CCT_REG_BITS[8] ), .A1N(N323), .B0(
        N303), .Y(A_AFTER_MUX[0]) );
  OAI221XLTF U337 ( .A0(N103), .A1(SCPU_CTRL_SPI_A_SPI[0]), .B0(N279), .B1(
        SCPU_CTRL_SPI_I_ADDR[0]), .C0(N270), .Y(N303) );
  AND2X2TF U338 ( .A(N323), .B(N93), .Y(N324) );
  NAND2X1TF U339 ( .A(\SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .B(N285), .Y(N219)
         );
  NOR2X2TF U340 ( .A(I_CTRL_BGN), .B(N103), .Y(N319) );
  INVX2TF U341 ( .A(N267), .Y(N423) );
  NOR2X1TF U342 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .B(N282), .Y(N335) );
  NAND3X1TF U343 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .B(
        \SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .C(N100), .Y(N353) );
  NAND2X1TF U344 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .B(N282), .Y(N337) );
  NOR2X1TF U345 ( .A(N392), .B(N290), .Y(SCPU_CTRL_SPI_PUT_N106) );
  AOI21X1TF U346 ( .A0(N429), .A1(N281), .B0(N284), .Y(N45) );
  OAI31X1TF U347 ( .A0(N346), .A1(N337), .A2(N339), .B0(N336), .Y(N212) );
  AOI32X1TF U348 ( .A0(N392), .A1(N100), .A2(N335), .B0(N289), .B1(N334), .Y(
        N336) );
  OAI21X1TF U349 ( .A0(N346), .A1(N345), .B0(N344), .Y(N209) );
  OAI21X1TF U350 ( .A0(N289), .A1(N394), .B0(\SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), 
        .Y(N344) );
  AOI211X1TF U351 ( .A0(N343), .A1(N289), .B0(N342), .C0(N273), .Y(N345) );
  AOI22X1TF U352 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .A1(N273), .B0(
        N427), .B1(N283), .Y(N33) );
  OAI32X1TF U353 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ), .A1(
        \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .A2(N427), .B0(N425), .B1(N278), 
        .Y(N36) );
  OAI32X1TF U354 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] ), .A1(N428), .A2(
        N427), .B0(N429), .B1(N281), .Y(N42) );
  NOR2X1TF U355 ( .A(N426), .B(N428), .Y(N429) );
  NOR2X1TF U356 ( .A(N100), .B(N346), .Y(N340) );
  AOI21X1TF U357 ( .A0(N289), .A1(N341), .B0(N392), .Y(N346) );
  NOR2X1TF U358 ( .A(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .B(N426), .Y(N425)
         );
  OAI211X1TF U359 ( .A0(N354), .A1(N292), .B0(N353), .C0(N352), .Y(N205) );
  AOI22X1TF U360 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ), .A1(N348), .B0(
        N349), .B1(N294), .Y(N208) );
  AOI21X1TF U361 ( .A0(N355), .A1(N338), .B0(N395), .Y(N348) );
  OAI211X1TF U362 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .A1(N352), .B0(
        N353), .C0(N351), .Y(N206) );
  OAI21X1TF U363 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .A1(N395), .B0(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .Y(N351) );
  INVX2TF U364 ( .A(N392), .Y(N394) );
  OAI31X1TF U365 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .A1(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .A2(N395), .B0(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ), .Y(N350) );
  NOR2X1TF U366 ( .A(N356), .B(N354), .Y(N395) );
  INVX2TF U367 ( .A(N347), .Y(N338) );
  NOR3X1TF U368 ( .A(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ), .B(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .C(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .Y(N347) );
  OAI22X1TF U369 ( .A0(I_CTRL_MODE[0]), .A1(N330), .B0(N329), .B1(N332), .Y(
        N215) );
  AOI21X1TF U370 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ), .A1(N328), .B0(
        N327), .Y(N329) );
  INVX2TF U371 ( .A(N332), .Y(N158) );
  NOR2X1TF U372 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .B(
        \SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .Y(N342) );
  AOI22X1TF U373 ( .A0(N296), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[1] ), .B0(N378), 
        .B1(I_CTRL_SO), .Y(N371) );
  AOI22X1TF U374 ( .A0(N296), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[4] ), .B0(N378), 
        .B1(\SCPU_CTRL_SPI_CCT_REG_BITS[3] ), .Y(N374) );
  AOI22X1TF U375 ( .A0(N296), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[8] ), .B0(N378), 
        .B1(\SCPU_CTRL_SPI_CCT_REG_BITS[7] ), .Y(N379) );
  AOI22X1TF U376 ( .A0(N296), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[7] ), .B0(N378), 
        .B1(\SCPU_CTRL_SPI_CCT_REG_BITS[6] ), .Y(N377) );
  AOI22X1TF U377 ( .A0(N296), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[2] ), .B0(N378), 
        .B1(\SCPU_CTRL_SPI_CCT_REG_BITS[1] ), .Y(N372) );
  AOI22X1TF U378 ( .A0(N296), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[5] ), .B0(N378), 
        .B1(\SCPU_CTRL_SPI_CCT_REG_BITS[4] ), .Y(N375) );
  AOI22X1TF U379 ( .A0(N296), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[3] ), .B0(N378), 
        .B1(\SCPU_CTRL_SPI_CCT_REG_BITS[2] ), .Y(N373) );
  AOI22X1TF U380 ( .A0(N296), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[6] ), .B0(N378), 
        .B1(\SCPU_CTRL_SPI_CCT_REG_BITS[5] ), .Y(N376) );
  NOR2X2TF U381 ( .A(N296), .B(N370), .Y(N378) );
  NAND2X2TF U382 ( .A(I_CTRL_BGN), .B(N370), .Y(N380) );
  NOR3X1TF U383 ( .A(I_CTRL_MODE[1]), .B(N369), .C(N219), .Y(N370) );
  NOR3X1TF U384 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ), .B(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ), .C(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .Y(N300) );
  NOR2X1TF U385 ( .A(N91), .B(\SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .Y(N220) );
  AOI32X1TF U386 ( .A0(N103), .A1(N270), .A2(SCPU_CTRL_SPI_D_WE), .B0(
        I_CTRL_BGN), .B1(N93), .Y(WEN_AFTER_MUX) );
  OAI32X1TF U387 ( .A0(N297), .A1(N333), .A2(N103), .B0(N426), .B1(N297), .Y(
        N213) );
  OAI31X1TF U388 ( .A0(SCPU_CTRL_SPI_A_SPI[3]), .A1(N422), .A2(N415), .B0(N414), .Y(N81) );
  AOI22X1TF U389 ( .A0(SCPU_CTRL_SPI_A_SPI[3]), .A1(N413), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[3] ), .B1(N298), .Y(N414) );
  AOI21X1TF U390 ( .A0(N273), .A1(N412), .B0(N298), .Y(N413) );
  OAI31X1TF U391 ( .A0(SCPU_CTRL_SPI_A_SPI[1]), .A1(N422), .A2(N293), .B0(N420), .Y(N79) );
  AOI22X1TF U392 ( .A0(SCPU_CTRL_SPI_A_SPI[1]), .A1(N419), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[1] ), .B1(N423), .Y(N420) );
  AOI21X1TF U393 ( .A0(N273), .A1(SCPU_CTRL_SPI_A_SPI[0]), .B0(N298), .Y(N419)
         );
  OAI31X1TF U394 ( .A0(SCPU_CTRL_SPI_A_SPI[6]), .A1(N422), .A2(N404), .B0(N403), .Y(N84) );
  AOI22X1TF U395 ( .A0(SCPU_CTRL_SPI_A_SPI[6]), .A1(N402), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[6] ), .B1(N423), .Y(N403) );
  AOI31X1TF U396 ( .A0(N273), .A1(N405), .A2(SCPU_CTRL_SPI_A_SPI[5]), .B0(N298), .Y(N402) );
  OAI31X1TF U397 ( .A0(SCPU_CTRL_SPI_A_SPI[5]), .A1(N422), .A2(N408), .B0(N407), .Y(N83) );
  AOI22X1TF U398 ( .A0(SCPU_CTRL_SPI_A_SPI[5]), .A1(N406), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[5] ), .B1(N423), .Y(N407) );
  AOI21X1TF U399 ( .A0(N273), .A1(N405), .B0(N298), .Y(N406) );
  OAI31X1TF U400 ( .A0(SCPU_CTRL_SPI_A_SPI[4]), .A1(N422), .A2(N411), .B0(N410), .Y(N82) );
  AOI22X1TF U401 ( .A0(SCPU_CTRL_SPI_A_SPI[4]), .A1(N409), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[4] ), .B1(N298), .Y(N410) );
  AOI31X1TF U402 ( .A0(N424), .A1(N412), .A2(SCPU_CTRL_SPI_A_SPI[3]), .B0(N298), .Y(N409) );
  OAI31X1TF U403 ( .A0(SCPU_CTRL_SPI_A_SPI[2]), .A1(N422), .A2(N418), .B0(N417), .Y(N80) );
  AOI22X1TF U404 ( .A0(SCPU_CTRL_SPI_A_SPI[2]), .A1(N416), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[2] ), .B1(N298), .Y(N417) );
  AOI31X1TF U405 ( .A0(N273), .A1(SCPU_CTRL_SPI_A_SPI[0]), .A2(
        SCPU_CTRL_SPI_A_SPI[1]), .B0(N298), .Y(N416) );
  OAI31X1TF U406 ( .A0(SCPU_CTRL_SPI_A_SPI[8]), .A1(N291), .A2(N399), .B0(N398), .Y(N86) );
  AOI22X1TF U407 ( .A0(SCPU_CTRL_SPI_A_SPI[8]), .A1(N397), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[8] ), .B1(N297), .Y(N398) );
  OAI21X1TF U408 ( .A0(SCPU_CTRL_SPI_A_SPI[7]), .A1(N422), .B0(N401), .Y(N397)
         );
  OAI21X1TF U409 ( .A0(N401), .A1(N291), .B0(N400), .Y(N85) );
  INVX2TF U410 ( .A(N415), .Y(N412) );
  OAI21X1TF U411 ( .A0(SCPU_CTRL_SPI_A_SPI[0]), .A1(N422), .B0(N421), .Y(N78)
         );
  INVX2TF U412 ( .A(N424), .Y(N427) );
  NAND2X2TF U413 ( .A(N424), .B(N267), .Y(N422) );
  INVX2TF U414 ( .A(N337), .Y(N333) );
  NOR2X1TF U415 ( .A(N383), .B(N389), .Y(SCPU_CTRL_SPI_I_DATAIN[1]) );
  NOR2X1TF U416 ( .A(N387), .B(N389), .Y(SCPU_CTRL_SPI_I_DATAIN[5]) );
  NOR2X1TF U417 ( .A(N382), .B(N389), .Y(SCPU_CTRL_SPI_I_DATAIN[0]) );
  NOR2X1TF U418 ( .A(N384), .B(N389), .Y(SCPU_CTRL_SPI_I_DATAIN[2]) );
  NOR2X1TF U419 ( .A(N386), .B(N389), .Y(SCPU_CTRL_SPI_I_DATAIN[4]) );
  NOR2X1TF U420 ( .A(N390), .B(N389), .Y(SCPU_CTRL_SPI_I_DATAIN[7]) );
  NOR2X1TF U421 ( .A(N388), .B(N389), .Y(SCPU_CTRL_SPI_I_DATAIN[6]) );
  NOR2X1TF U422 ( .A(N385), .B(N389), .Y(SCPU_CTRL_SPI_I_DATAIN[3]) );
  INVX2TF U423 ( .A(Q_FROM_SRAM[7]), .Y(N390) );
  AOI22X1TF U424 ( .A0(N320), .A1(SCPU_CTRL_SPI_D_ADDR[8]), .B0(N323), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[16] ), .Y(N321) );
  AOI22X1TF U425 ( .A0(SCPU_CTRL_SPI_A_SPI[8]), .A1(N319), .B0(N318), .B1(
        SCPU_CTRL_SPI_I_ADDR[8]), .Y(N322) );
  AOI22X1TF U426 ( .A0(N320), .A1(SCPU_CTRL_SPI_D_ADDR[7]), .B0(N323), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[15] ), .Y(N316) );
  AOI22X1TF U427 ( .A0(SCPU_CTRL_SPI_A_SPI[7]), .A1(N319), .B0(N318), .B1(
        SCPU_CTRL_SPI_I_ADDR[7]), .Y(N317) );
  AOI22X1TF U428 ( .A0(N320), .A1(SCPU_CTRL_SPI_D_ADDR[6]), .B0(N323), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[14] ), .Y(N314) );
  AOI22X1TF U429 ( .A0(SCPU_CTRL_SPI_A_SPI[6]), .A1(N319), .B0(N318), .B1(
        SCPU_CTRL_SPI_I_ADDR[6]), .Y(N315) );
  AOI22X1TF U430 ( .A0(N320), .A1(SCPU_CTRL_SPI_D_ADDR[5]), .B0(N323), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[13] ), .Y(N312) );
  AOI22X1TF U431 ( .A0(SCPU_CTRL_SPI_A_SPI[5]), .A1(N319), .B0(N318), .B1(
        SCPU_CTRL_SPI_I_ADDR[5]), .Y(N313) );
  AOI22X1TF U432 ( .A0(N320), .A1(SCPU_CTRL_SPI_D_ADDR[4]), .B0(N323), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[12] ), .Y(N310) );
  AOI22X1TF U433 ( .A0(SCPU_CTRL_SPI_A_SPI[4]), .A1(N319), .B0(N318), .B1(
        SCPU_CTRL_SPI_I_ADDR[4]), .Y(N311) );
  AOI22X1TF U434 ( .A0(N320), .A1(SCPU_CTRL_SPI_D_ADDR[3]), .B0(N323), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[11] ), .Y(N308) );
  AOI22X1TF U435 ( .A0(SCPU_CTRL_SPI_A_SPI[3]), .A1(N319), .B0(N318), .B1(
        SCPU_CTRL_SPI_I_ADDR[3]), .Y(N309) );
  AOI22X1TF U436 ( .A0(N320), .A1(SCPU_CTRL_SPI_D_ADDR[2]), .B0(N323), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[10] ), .Y(N306) );
  AOI22X1TF U437 ( .A0(SCPU_CTRL_SPI_A_SPI[2]), .A1(N319), .B0(N318), .B1(
        SCPU_CTRL_SPI_I_ADDR[2]), .Y(N307) );
  AOI22X1TF U438 ( .A0(N320), .A1(SCPU_CTRL_SPI_D_ADDR[1]), .B0(N323), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[9] ), .Y(N304) );
  AOI22X1TF U439 ( .A0(SCPU_CTRL_SPI_A_SPI[1]), .A1(N319), .B0(N318), .B1(
        SCPU_CTRL_SPI_I_ADDR[1]), .Y(N305) );
  OAI21X1TF U440 ( .A0(N388), .A1(N367), .B0(N363), .Y(N198) );
  AOI22X1TF U441 ( .A0(N365), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[6]), .B0(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[7]), .B1(N364), .Y(N363) );
  INVX2TF U442 ( .A(Q_FROM_SRAM[6]), .Y(N388) );
  OAI21X1TF U443 ( .A0(N382), .A1(N367), .B0(N366), .Y(N197) );
  AOI22X1TF U444 ( .A0(N365), .A1(I_SPI_SO), .B0(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[1]), .B1(N364), .Y(N366) );
  INVX2TF U445 ( .A(Q_FROM_SRAM[0]), .Y(N382) );
  OAI21X1TF U446 ( .A0(N386), .A1(N367), .B0(N361), .Y(N200) );
  AOI22X1TF U447 ( .A0(N365), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[4]), .B0(N364), 
        .B1(SCPU_CTRL_SPI_PUT_SRAM_REGS[5]), .Y(N361) );
  INVX2TF U448 ( .A(Q_FROM_SRAM[4]), .Y(N386) );
  OAI21X1TF U449 ( .A0(N385), .A1(N367), .B0(N360), .Y(N201) );
  AOI22X1TF U450 ( .A0(N365), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[3]), .B0(N364), 
        .B1(SCPU_CTRL_SPI_PUT_SRAM_REGS[4]), .Y(N360) );
  INVX2TF U451 ( .A(Q_FROM_SRAM[3]), .Y(N385) );
  OAI21X1TF U452 ( .A0(N383), .A1(N367), .B0(N358), .Y(N203) );
  AOI22X1TF U453 ( .A0(N365), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[1]), .B0(N364), 
        .B1(SCPU_CTRL_SPI_PUT_SRAM_REGS[2]), .Y(N358) );
  INVX2TF U454 ( .A(Q_FROM_SRAM[1]), .Y(N383) );
  OAI21X1TF U455 ( .A0(N387), .A1(N367), .B0(N362), .Y(N199) );
  AOI22X1TF U456 ( .A0(N365), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[5]), .B0(N364), 
        .B1(SCPU_CTRL_SPI_PUT_SRAM_REGS[6]), .Y(N362) );
  INVX2TF U457 ( .A(Q_FROM_SRAM[5]), .Y(N387) );
  OAI21X1TF U458 ( .A0(N384), .A1(N367), .B0(N359), .Y(N202) );
  AOI22X1TF U459 ( .A0(N365), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[2]), .B0(N364), 
        .B1(SCPU_CTRL_SPI_PUT_SRAM_REGS[3]), .Y(N359) );
  NOR2X2TF U460 ( .A(N297), .B(N357), .Y(N364) );
  INVX2TF U461 ( .A(N355), .Y(N357) );
  INVX2TF U462 ( .A(N335), .Y(N341) );
  NAND3X2TF U463 ( .A(N269), .B(N267), .C(N356), .Y(N367) );
  INVX2TF U464 ( .A(N353), .Y(N356) );
  INVX2TF U465 ( .A(Q_FROM_SRAM[2]), .Y(N384) );
  NOR2X1TF U466 ( .A(N100), .B(N337), .Y(N221) );
  NOR3X1TF U467 ( .A(N102), .B(N103), .C(N286), .Y(I_SCLK1) );
  NOR3X1TF U468 ( .A(\SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .B(N102), .C(N103), 
        .Y(I_SCLK2) );
  INVX2TF U469 ( .A(N272), .Y(N391) );
  CLKBUFX2TF U470 ( .A(N297), .Y(N298) );
  OAI2BB1X1TF U471 ( .A0N(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .A1N(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ), .B0(N299), .Y(
        SCPU_CTRL_SPI_CCT_N49) );
  NOR2BX1TF U472 ( .AN(SCPU_CTRL_SPI_CEN), .B(N270), .Y(CEN_AFTER_MUX) );
  AO22X1TF U473 ( .A0(N324), .A1(I_CTRL_SO), .B0(SCPU_CTRL_SPI_D_DATAOUT[0]), 
        .B1(N270), .Y(D_AFTER_MUX[0]) );
  AO22X1TF U474 ( .A0(N324), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[1] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[1]), .B1(N270), .Y(D_AFTER_MUX[1]) );
  AO22X1TF U475 ( .A0(N324), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[2] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[2]), .B1(N270), .Y(D_AFTER_MUX[2]) );
  AO22X1TF U476 ( .A0(N324), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[3] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[3]), .B1(N269), .Y(D_AFTER_MUX[3]) );
  AO22X1TF U477 ( .A0(N324), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[4] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[4]), .B1(N270), .Y(D_AFTER_MUX[4]) );
  AO22X1TF U478 ( .A0(N324), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[5] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[5]), .B1(N269), .Y(D_AFTER_MUX[5]) );
  AO22X1TF U479 ( .A0(N324), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[6] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[6]), .B1(N270), .Y(D_AFTER_MUX[6]) );
  AO22X1TF U480 ( .A0(N324), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[7] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[7]), .B1(N270), .Y(D_AFTER_MUX[7]) );
  NAND2BX1TF U481 ( .AN(N219), .B(I_CTRL_MODE[1]), .Y(N218) );
  OAI221XLTF U482 ( .A0(\SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .A1(I_LOAD_N), 
        .B0(N368), .B1(N369), .C0(I_CTRL_BGN), .Y(N325) );
  NAND3BX1TF U483 ( .AN(I_LOAD_N), .B(N302), .C(N326), .Y(N330) );
  AO21X1TF U484 ( .A0(I_CTRL_MODE[0]), .A1(I_CTRL_MODE[1]), .B0(N330), .Y(N331) );
  NAND3X1TF U485 ( .A(N280), .B(N283), .C(N278), .Y(N428) );
  NAND3BX1TF U486 ( .AN(N428), .B(N281), .C(N284), .Y(N339) );
  OAI222X1TF U487 ( .A0(N427), .A1(N346), .B0(N341), .B1(N343), .C0(N282), 
        .C1(N340), .Y(N210) );
  NAND2X1TF U488 ( .A(N347), .B(N354), .Y(N349) );
  NAND3X1TF U489 ( .A(N353), .B(N350), .C(N349), .Y(N207) );
  NAND2X1TF U490 ( .A(N354), .B(N292), .Y(N352) );
  OAI2BB2XLTF U491 ( .B0(N390), .B1(N367), .A0N(N365), .A1N(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[7]), .Y(N204) );
  AO22X1TF U492 ( .A0(N272), .A1(SCPU_CTRL_SPI_FOUT[0]), .B0(N295), .B1(
        I_ADC_PI[0]), .Y(SCPU_CTRL_SPI_IO_DATAINA[0]) );
  AO22X1TF U493 ( .A0(N272), .A1(SCPU_CTRL_SPI_FOUT[10]), .B0(N391), .B1(
        I_ADC_PI[10]), .Y(SCPU_CTRL_SPI_IO_DATAINA[10]) );
  AO22X1TF U494 ( .A0(N272), .A1(SCPU_CTRL_SPI_FOUT[11]), .B0(N391), .B1(
        I_ADC_PI[11]), .Y(SCPU_CTRL_SPI_IO_DATAINA[11]) );
  AO22X1TF U495 ( .A0(N271), .A1(SCPU_CTRL_SPI_FOUT[12]), .B0(N295), .B1(
        I_ADC_PI[12]), .Y(SCPU_CTRL_SPI_IO_DATAINA[12]) );
  NOR2BX1TF U496 ( .AN(I_ADC_PI[13]), .B(N271), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[13]) );
  NOR2BX1TF U497 ( .AN(I_ADC_PI[14]), .B(N272), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[14]) );
  NOR2BX1TF U498 ( .AN(I_ADC_PI[15]), .B(N271), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[15]) );
  AO22X1TF U499 ( .A0(N271), .A1(SCPU_CTRL_SPI_FOUT[1]), .B0(N391), .B1(
        I_ADC_PI[1]), .Y(SCPU_CTRL_SPI_IO_DATAINA[1]) );
  AO22X1TF U500 ( .A0(N271), .A1(SCPU_CTRL_SPI_FOUT[2]), .B0(N391), .B1(
        I_ADC_PI[2]), .Y(SCPU_CTRL_SPI_IO_DATAINA[2]) );
  AO22X1TF U501 ( .A0(N272), .A1(SCPU_CTRL_SPI_FOUT[3]), .B0(N295), .B1(
        I_ADC_PI[3]), .Y(SCPU_CTRL_SPI_IO_DATAINA[3]) );
  AO22X1TF U502 ( .A0(N271), .A1(SCPU_CTRL_SPI_FOUT[4]), .B0(N391), .B1(
        I_ADC_PI[4]), .Y(SCPU_CTRL_SPI_IO_DATAINA[4]) );
  AO22X1TF U503 ( .A0(N272), .A1(SCPU_CTRL_SPI_FOUT[5]), .B0(N391), .B1(
        I_ADC_PI[5]), .Y(SCPU_CTRL_SPI_IO_DATAINA[5]) );
  AO22X1TF U504 ( .A0(N271), .A1(SCPU_CTRL_SPI_FOUT[6]), .B0(N391), .B1(
        I_ADC_PI[6]), .Y(SCPU_CTRL_SPI_IO_DATAINA[6]) );
  AO22X1TF U505 ( .A0(N272), .A1(SCPU_CTRL_SPI_FOUT[7]), .B0(N391), .B1(
        I_ADC_PI[7]), .Y(SCPU_CTRL_SPI_IO_DATAINA[7]) );
  AO22X1TF U506 ( .A0(N271), .A1(SCPU_CTRL_SPI_FOUT[8]), .B0(N391), .B1(
        I_ADC_PI[8]), .Y(SCPU_CTRL_SPI_IO_DATAINA[8]) );
  AO22X1TF U507 ( .A0(N272), .A1(SCPU_CTRL_SPI_FOUT[9]), .B0(N391), .B1(
        I_ADC_PI[9]), .Y(SCPU_CTRL_SPI_IO_DATAINA[9]) );
  OAI2BB2XLTF U508 ( .B0(N286), .B1(N102), .A0N(N286), .A1N(
        SCPU_CTRL_SPI_PUT_N106), .Y(SCPU_CTRL_SPI_PUT_N107) );
  NAND2X1TF U509 ( .A(N102), .B(N286), .Y(N393) );
  NAND3X1TF U510 ( .A(SCPU_CTRL_SPI_A_SPI[2]), .B(SCPU_CTRL_SPI_A_SPI[0]), .C(
        SCPU_CTRL_SPI_A_SPI[1]), .Y(N415) );
  NAND2X1TF U511 ( .A(N412), .B(SCPU_CTRL_SPI_A_SPI[3]), .Y(N411) );
  NOR2BX1TF U512 ( .AN(SCPU_CTRL_SPI_A_SPI[4]), .B(N411), .Y(N405) );
  NAND2X1TF U513 ( .A(N405), .B(SCPU_CTRL_SPI_A_SPI[5]), .Y(N404) );
  NOR2BX1TF U514 ( .AN(SCPU_CTRL_SPI_A_SPI[6]), .B(N404), .Y(N396) );
  NAND2BX1TF U515 ( .AN(N422), .B(N396), .Y(N399) );
  OAI2BB1X1TF U516 ( .A0N(N424), .A1N(N396), .B0(N267), .Y(N401) );
  AOI2BB2X1TF U517 ( .B0(\SCPU_CTRL_SPI_IO_DATAOUTA[7] ), .B1(N297), .A0N(
        SCPU_CTRL_SPI_A_SPI[7]), .A1N(N399), .Y(N400) );
  NAND2X1TF U519 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[3] ), .B(N423), .Y(N41) );
  NAND2X1TF U520 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[2] ), .B(N297), .Y(N38) );
  NAND2X1TF U521 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[1] ), .B(N297), .Y(N35) );
  NAND2X1TF U522 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[0] ), .B(N298), .Y(N32) );
endmodule

