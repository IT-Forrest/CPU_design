
module SHARE_SUPERALU_VG ( CLK, RST_N, X_IN, Y_IN, ALU_START, ALU_TYPE, MODE_TYPE, 
        OFFSET, FOUT, POUT, ALU_IS_DONE );
  input [12:0] X_IN;
  input [12:0] Y_IN;
  input [2:0] ALU_TYPE;
  input [1:0] MODE_TYPE;
  input [9:0] OFFSET;
  output [12:0] FOUT;
  output [12:0] POUT;
  input CLK, RST_N, ALU_START;
  output ALU_IS_DONE;
  wire   POST_WORK, PRE_WORK, \INDEX[2] , \RSHT_BITS[3] , SIGN_Y, C152_DATA4_0,
         C152_DATA4_1, C152_DATA4_2, C152_DATA4_3, C152_DATA4_4, C152_DATA4_5,
         C152_DATA4_6, C152_DATA4_7, C152_DATA4_8, C152_DATA4_9, C152_DATA4_10,
         C152_DATA4_11, N73, N74, N90, N91, N92, N121, N122, N123, N124, N128,
         N129, N657, N658, N659, N660, N661, N662, N663, N664, N665, N666,
         N667, N668, N669, N670, N671, N672, N673, N674, N675, N676, N677,
         N678, N679, N680, N681, N682, N683, N684, N685, N686, N687, N688,
         N689, N690, N691, N692, N693, N694, N695, N696, N697, N698, N699,
         N700, N701, N702, N703, N704, N705, N706, N707, N708, N709, N710,
         N711, N712, N713, N714, N715, N716, N717, N718, N719, N720, N721,
         N722, N723, N724, N725, N726, C2_Z_11, C2_Z_10, C2_Z_9, C2_Z_8,
         C2_Z_7, C2_Z_6, C2_Z_5, C2_Z_4, C2_Z_3, C2_Z_2, C2_Z_1,
         DP_OP_333_124_4748_N57, DP_OP_333_124_4748_N43,
         DP_OP_333_124_4748_N28, DP_OP_333_124_4748_N27,
         DP_OP_333_124_4748_N26, DP_OP_333_124_4748_N25,
         DP_OP_333_124_4748_N24, DP_OP_333_124_4748_N23,
         DP_OP_333_124_4748_N22, DP_OP_333_124_4748_N21,
         DP_OP_333_124_4748_N20, DP_OP_333_124_4748_N19,
         DP_OP_333_124_4748_N18, DP_OP_333_124_4748_N12,
         DP_OP_333_124_4748_N11, DP_OP_333_124_4748_N10, DP_OP_333_124_4748_N9,
         DP_OP_333_124_4748_N8, DP_OP_333_124_4748_N7, DP_OP_333_124_4748_N6,
         DP_OP_333_124_4748_N5, DP_OP_333_124_4748_N4, DP_OP_333_124_4748_N3,
         DP_OP_333_124_4748_N2, DP_OP_333_124_4748_N1, INTADD_0_CI,
         \INTADD_0_SUM[6] , \INTADD_0_SUM[5] , \INTADD_0_SUM[4] ,
         \INTADD_0_SUM[3] , \INTADD_0_SUM[2] , \INTADD_0_SUM[1] ,
         \INTADD_0_SUM[0] , INTADD_0_N7, INTADD_0_N6, INTADD_0_N5, INTADD_0_N4,
         INTADD_0_N3, INTADD_0_N2, INTADD_0_N1, ADD_X_132_1_N13,
         ADD_X_132_1_N12, ADD_X_132_1_N11, ADD_X_132_1_N10, ADD_X_132_1_N9,
         ADD_X_132_1_N8, ADD_X_132_1_N7, ADD_X_132_1_N6, ADD_X_132_1_N5,
         ADD_X_132_1_N4, ADD_X_132_1_N3, ADD_X_132_1_N2, N1, N2, N3, N4, N5,
         N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20,
         N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32, N33, N34,
         N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48,
         N49, N50, N51, N52, N53, N54, N55, N56, N78, N79, N80, N81, N82, N83,
         N84, N85, N86, N87, N88, N89, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N114, N115, N116, N117, N118, N119, N120, N125, N126,
         N127, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139,
         N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161,
         N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172,
         N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183,
         N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194,
         N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205,
         N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216,
         N217, N218, N219, N220, N221, N222, N223, N224, N225, N226, N227,
         N228, N229, N230, N231, N232, N233, N234, N235, N236, N237, N238,
         N239, N240, N241, N242, N243, N244, N245, N246, N247, N248, N249,
         N250, N251, N252, N253, N254, N255, N256, N257, N258, N259, N260,
         N261, N262, N263, N264, N265, N266, N267, N268, N269, N270, N271,
         N272, N273, N274, N275, N276, N277, N278, N279, N280, N281, N282,
         N283, N284, N285, N286, N287, N288, N289, N290, N291, N292, N293,
         N294, N295, N296, N297, N298, N299, N300, N301, N302, N303, N304,
         N305, N306, N307, N308, N309, N310, N311, N312, N313, N314, N315,
         N316, N317, N318, N319, N320, N321, N322, N323, N324, N325, N326,
         N327, N328, N329, N330, N331, N332, N333, N334, N335, N336, N337,
         N338, N339, N340, N341, N342, N343, N344, N345, N346, N347, N348,
         N349, N350, N351, N352, N353, N354, N355, N356, N357, N358, N359,
         N360, N361, N362, N363, N364, N365, N366, N367, N368, N369, N370,
         N371, N372, N373, N374, N375, N376, N377, N378, N379, N380, N381,
         N382, N383, N384, N385, N386, N387, N388, N389, N390, N391, N392,
         N393, N394, N395, N396, N397, N398, N399, N400, N401, N402, N403,
         N404, N405, N406, N407, N408, N409, N410, N411, N412, N413, N414,
         N415, N416, N417, N418, N419, N420, N421, N422, N423, N424, N425,
         N426, N427, N428, N429, N430, N431, N432, N433, N434, N435, N436,
         N437, N438, N439, N440, N441, N442, N443, N444, N445, N446, N447,
         N448, N449, N450, N451, N452, N453, N454, N455, N456, N457, N458,
         N459, N460, N461, N462, N463, N464, N465, N466, N467, N468, N469,
         N470, N471, N472, N473, N474, N475, N476, N477, N478, N479, N480,
         N481, N482, N483, N484, N485, N486, N487, N488, N489, N490, N491,
         N492, N493, N494, N495, N496, N497, N498, N499, N500, N501, N502,
         N503, N504, N505, N506, N507, N508, N509, N510, N511, N512, N513,
         N514, N515, N516, N517, N518, N519, N520, N521, N522, N523, N524,
         N525, N526, N527, N528, N529, N530, N531, N532, N533, N534, N535,
         N536, N537, N538, N539, N540, N541, N542, N543, N544, N545, N546,
         N547, N548, N549, N550, N551, N552, N553, N554, N555, N556, N557,
         N558, N559, N560, N561, N562, N563, N564, N565, N566, N567, N568,
         N569, N570, N571, N572, N573, N574, N575, N576, N577, N578, N579,
         N580, N581, N582, N583, N584, N585, N586, N587, N588, N589, N590,
         N591, N592, N593, N594, N595, N596, N597, N598, N599, N600, N601,
         N602, N603, N604, N605, N606, N607, N608, N609, N610, N611, N612,
         N613, N614, N615, N616, N617, N618, N619, N620, N621, N622, N623,
         N624, N625, N626, N627, N628, N629, N630, N631, N632, N633, N634,
         N635, N636, N637, N638, N639, N640, N641, N642, N643, N644, N645,
         N646, N647, N648, N649, N650, N651, N652, N653, N654, N655, N656,
         N727, N728, N729, N730, N731, N732, N733, N734, N735, N736, N737,
         N738, N739, N740, N741, N742, N743, N744, N745, N746, N747, N748,
         N749, N750, N751, N752, N753, N754, N755, N756, N757, N758, N759,
         N760, N761, N762, N763, N764, N765, N766, N767, N768, N769, N770,
         N771, N772, N773, N774, N775, N776, N777, N778, N779, N780, N781,
         N782, N783, N784, N785, N786, N787, N788, N789, N790, N791, N792,
         N793, N794, N795, N796, N797, N798, N799, N800, N801, N802, N803,
         N804, N805, N806, N807, N808, N809, N810, N811, N812, N813, N814,
         N815, N816, N817, N818, N819, N820, N821, N822, N823, N824, N825,
         N826, N827, N828, N829, N830, N831, N832, N833, N834, N835, N836,
         N837, N838, N839, N840, N841, N842, N843, N844, N845, N846, N847,
         N848, N849, N850, N851, N852, N853, N854, N855, N856, N857, N858,
         N859, N860, N861, N862, N863, N864, N865, N866, N867, N868, N869,
         N870, N871, N872, N873, N874, N875, N876, N877, N878, N879, N880,
         N881, N882, N883, N884, N885, N886, N887, N888, N889, N890, N891,
         N892, N893, N894, N895, N896, N897, N898, N899, N900, N901, N902,
         N903, N904, N905, N906, N907, N908, N909, N910, N911, N912, N913,
         N914, N915, N916, N917, N918, N919, N920, N921, N922, N923, N924,
         N925, N926, N927, N928, N929, N930, N931, N932, N933, N934, N935,
         N936, N937, N938, N939, N940, N941, N942, N943, N944, N945, N946,
         N947, N948, N949, N950, N951, N952, N953, N954, N955, N956, N957,
         N958, N959, N960, N961, N962, N963, N964, N965, N966, N967, N968,
         N969, N970, N971, N972, N973, N974, N975, N976, N977, N978, N979,
         N980, N981, N982, N983, N984, N985, N986, N987, N988, N989, N990,
         N991, N992, N993, N994, N995, N996, N997, N998, N999, N1000, N1001,
         N1002, N1003, N1004, N1005, N1006, N1007, N1008, N1009, N1010, N1011,
         N1012, N1013, N1014, N1015, N1016, N1017, N1018, N1019;
  wire   [12:9] XTEMP;
  wire   [12:0] DIVISION_HEAD;
  wire   [8:0] DIVISION_REMA;
  wire   [12:0] OPER_A;
  wire   [12:0] OPER_B;
  wire   [12:0] SUM_AB;
  wire   [12:0] ZTEMP;
  wire   [3:2] STEP;

  XOR2X1TF \DP_OP_333_124_4748/U27  ( .A(N78), .B(C2_Z_1), .Y(
        DP_OP_333_124_4748_N28) );
  XOR2X1TF \DP_OP_333_124_4748/U26  ( .A(N78), .B(C2_Z_2), .Y(
        DP_OP_333_124_4748_N27) );
  XOR2X1TF \DP_OP_333_124_4748/U25  ( .A(N78), .B(C2_Z_3), .Y(
        DP_OP_333_124_4748_N26) );
  XOR2X1TF \DP_OP_333_124_4748/U24  ( .A(N125), .B(C2_Z_4), .Y(
        DP_OP_333_124_4748_N25) );
  XOR2X1TF \DP_OP_333_124_4748/U23  ( .A(N78), .B(C2_Z_5), .Y(
        DP_OP_333_124_4748_N24) );
  XOR2X1TF \DP_OP_333_124_4748/U22  ( .A(N125), .B(C2_Z_6), .Y(
        DP_OP_333_124_4748_N23) );
  XOR2X1TF \DP_OP_333_124_4748/U21  ( .A(N78), .B(C2_Z_7), .Y(
        DP_OP_333_124_4748_N22) );
  XOR2X1TF \DP_OP_333_124_4748/U20  ( .A(N125), .B(C2_Z_8), .Y(
        DP_OP_333_124_4748_N21) );
  XOR2X1TF \DP_OP_333_124_4748/U19  ( .A(N78), .B(C2_Z_9), .Y(
        DP_OP_333_124_4748_N20) );
  XOR2X1TF \DP_OP_333_124_4748/U18  ( .A(N125), .B(C2_Z_10), .Y(
        DP_OP_333_124_4748_N19) );
  XOR2X1TF \DP_OP_333_124_4748/U17  ( .A(N78), .B(C2_Z_11), .Y(
        DP_OP_333_124_4748_N18) );
  ADDHXLTF \DP_OP_333_124_4748/U12  ( .A(DP_OP_333_124_4748_N28), .B(
        DP_OP_333_124_4748_N12), .CO(DP_OP_333_124_4748_N11), .S(C152_DATA4_1)
         );
  ADDHXLTF \DP_OP_333_124_4748/U11  ( .A(DP_OP_333_124_4748_N27), .B(
        DP_OP_333_124_4748_N11), .CO(DP_OP_333_124_4748_N10), .S(C152_DATA4_2)
         );
  ADDHXLTF \DP_OP_333_124_4748/U10  ( .A(DP_OP_333_124_4748_N26), .B(
        DP_OP_333_124_4748_N10), .CO(DP_OP_333_124_4748_N9), .S(C152_DATA4_3)
         );
  ADDHXLTF \DP_OP_333_124_4748/U9  ( .A(DP_OP_333_124_4748_N25), .B(
        DP_OP_333_124_4748_N9), .CO(DP_OP_333_124_4748_N8), .S(C152_DATA4_4)
         );
  ADDHXLTF \DP_OP_333_124_4748/U8  ( .A(DP_OP_333_124_4748_N24), .B(
        DP_OP_333_124_4748_N8), .CO(DP_OP_333_124_4748_N7), .S(C152_DATA4_5)
         );
  ADDHXLTF \DP_OP_333_124_4748/U7  ( .A(DP_OP_333_124_4748_N23), .B(
        DP_OP_333_124_4748_N7), .CO(DP_OP_333_124_4748_N6), .S(C152_DATA4_6)
         );
  ADDHXLTF \DP_OP_333_124_4748/U6  ( .A(DP_OP_333_124_4748_N22), .B(
        DP_OP_333_124_4748_N6), .CO(DP_OP_333_124_4748_N5), .S(C152_DATA4_7)
         );
  ADDHXLTF \DP_OP_333_124_4748/U5  ( .A(DP_OP_333_124_4748_N21), .B(
        DP_OP_333_124_4748_N5), .CO(DP_OP_333_124_4748_N4), .S(C152_DATA4_8)
         );
  ADDHXLTF \DP_OP_333_124_4748/U4  ( .A(DP_OP_333_124_4748_N20), .B(
        DP_OP_333_124_4748_N4), .CO(DP_OP_333_124_4748_N3), .S(C152_DATA4_9)
         );
  ADDHXLTF \DP_OP_333_124_4748/U3  ( .A(DP_OP_333_124_4748_N19), .B(
        DP_OP_333_124_4748_N3), .CO(DP_OP_333_124_4748_N2), .S(C152_DATA4_10)
         );
  ADDHXLTF \DP_OP_333_124_4748/U2  ( .A(DP_OP_333_124_4748_N18), .B(
        DP_OP_333_124_4748_N2), .CO(DP_OP_333_124_4748_N1), .S(C152_DATA4_11)
         );
  CMPR32X2TF \intadd_0/U8  ( .A(X_IN[1]), .B(DIVISION_HEAD[5]), .C(INTADD_0_CI), .CO(INTADD_0_N7), .S(\INTADD_0_SUM[0] ) );
  CMPR32X2TF \intadd_0/U7  ( .A(X_IN[2]), .B(DIVISION_HEAD[6]), .C(INTADD_0_N7), .CO(INTADD_0_N6), .S(\INTADD_0_SUM[1] ) );
  CMPR32X2TF \intadd_0/U6  ( .A(X_IN[3]), .B(DIVISION_HEAD[7]), .C(INTADD_0_N6), .CO(INTADD_0_N5), .S(\INTADD_0_SUM[2] ) );
  CMPR32X2TF \intadd_0/U5  ( .A(X_IN[4]), .B(DIVISION_HEAD[8]), .C(INTADD_0_N5), .CO(INTADD_0_N4), .S(\INTADD_0_SUM[3] ) );
  CMPR32X2TF \intadd_0/U4  ( .A(X_IN[5]), .B(DIVISION_HEAD[9]), .C(INTADD_0_N4), .CO(INTADD_0_N3), .S(\INTADD_0_SUM[4] ) );
  CMPR32X2TF \intadd_0/U3  ( .A(X_IN[6]), .B(DIVISION_HEAD[10]), .C(
        INTADD_0_N3), .CO(INTADD_0_N2), .S(\INTADD_0_SUM[5] ) );
  CMPR32X2TF \intadd_0/U2  ( .A(X_IN[7]), .B(DIVISION_HEAD[11]), .C(
        INTADD_0_N2), .CO(INTADD_0_N1), .S(\INTADD_0_SUM[6] ) );
  DFFRX2TF \rsht_bits_reg[3]  ( .D(N704), .CK(CLK), .RN(RST_N), .Q(
        \RSHT_BITS[3] ), .QN(N189) );
  DFFRX2TF \wtemp_reg[9]  ( .D(N673), .CK(CLK), .RN(RST_N), .Q(OPER_B[9]), 
        .QN(N188) );
  DFFRX2TF \wtemp_reg[12]  ( .D(N724), .CK(CLK), .RN(RST_N), .Q(OPER_B[12]), 
        .QN(N187) );
  DFFRX2TF \index_reg[3]  ( .D(N725), .CK(CLK), .RN(RST_N), .Q(N186), .QN(N124) );
  DFFRX2TF \wtemp_reg[11]  ( .D(N671), .CK(CLK), .RN(RST_N), .Q(OPER_B[11]), 
        .QN(N185) );
  DFFRX2TF \wtemp_reg[0]  ( .D(N682), .CK(CLK), .RN(RST_N), .Q(OPER_B[0]), 
        .QN(N184) );
  DFFRX2TF \wtemp_reg[3]  ( .D(N679), .CK(CLK), .RN(RST_N), .Q(OPER_B[3]), 
        .QN(N183) );
  DFFRX2TF \wtemp_reg[1]  ( .D(N681), .CK(CLK), .RN(RST_N), .Q(OPER_B[1]), 
        .QN(N182) );
  DFFRX2TF \index_reg[1]  ( .D(N699), .CK(CLK), .RN(RST_N), .Q(N181), .QN(N128) );
  DFFRX2TF \rsht_bits_reg[0]  ( .D(N703), .CK(CLK), .RN(RST_N), .Q(N180), .QN(
        N92) );
  DFFRX2TF \ytemp_reg[0]  ( .D(N705), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[0]), .QN(N179) );
  DFFRX2TF sign_y_reg ( .D(N694), .CK(CLK), .RN(RST_N), .Q(SIGN_Y), .QN(N178)
         );
  DFFRX2TF \wtemp_reg[4]  ( .D(N678), .CK(CLK), .RN(RST_N), .Q(OPER_B[4]), 
        .QN(N177) );
  DFFRX2TF \xtemp_reg[8]  ( .D(N711), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[12]), .QN(N176) );
  DFFSX2TF pre_work_reg ( .D(N695), .CK(CLK), .SN(RST_N), .Q(PRE_WORK), .QN(
        N175) );
  DFFRX2TF \ytemp_reg[6]  ( .D(N688), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[6]), .QN(N174) );
  DFFRX2TF \ytemp_reg[10]  ( .D(N684), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[1]), .QN(N173) );
  DFFRX2TF \ytemp_reg[2]  ( .D(N692), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[2]), .QN(N172) );
  DFFRX2TF \xtemp_reg[12]  ( .D(N723), .CK(CLK), .RN(RST_N), .Q(XTEMP[12]), 
        .QN(N171) );
  DFFRX2TF \ytemp_reg[4]  ( .D(N690), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[4]), .QN(N170) );
  DFFRX2TF \ytemp_reg[9]  ( .D(N685), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[0]), .QN(N169) );
  DFFRX2TF \ytemp_reg[7]  ( .D(N687), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[7]), .QN(N168) );
  DFFRX2TF \ytemp_reg[5]  ( .D(N689), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[5]), .QN(N167) );
  DFFRX2TF \ytemp_reg[3]  ( .D(N691), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[3]), .QN(N166) );
  DFFRX2TF \step_reg[0]  ( .D(N697), .CK(CLK), .RN(RST_N), .Q(N165), .QN(N122)
         );
  DFFRX2TF \ytemp_reg[11]  ( .D(N683), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[2]), .QN(N163) );
  DFFRX2TF SEL_SRC_reg ( .D(N720), .CK(CLK), .RN(RST_N), .Q(POST_WORK), .QN(
        N162) );
  DFFRX2TF \wtemp_reg[10]  ( .D(N672), .CK(CLK), .RN(RST_N), .Q(OPER_B[10]), 
        .QN(N161) );
  DFFRX2TF \wtemp_reg[8]  ( .D(N674), .CK(CLK), .RN(RST_N), .Q(OPER_B[8]), 
        .QN(N160) );
  DFFRX2TF \ytemp_reg[1]  ( .D(N693), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[1]), .QN(N159) );
  DFFRX2TF \rsht_bits_reg[1]  ( .D(N702), .CK(CLK), .RN(RST_N), .Q(N158), .QN(
        N91) );
  DFFRX2TF \index_reg[0]  ( .D(N726), .CK(CLK), .RN(RST_N), .Q(N157), .QN(N129) );
  DFFRX2TF \wtemp_reg[2]  ( .D(N680), .CK(CLK), .RN(RST_N), .Q(OPER_B[2]), 
        .QN(N156) );
  DFFRX2TF \xtemp_reg[11]  ( .D(N708), .CK(CLK), .RN(RST_N), .Q(XTEMP[11]), 
        .QN(N155) );
  DFFRX2TF \xtemp_reg[6]  ( .D(N713), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[10]), .QN(N154) );
  DFFRX2TF \xtemp_reg[0]  ( .D(N719), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[4]), .QN(N153) );
  DFFRX2TF \xtemp_reg[2]  ( .D(N717), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[6]), .QN(N152) );
  DFFRX2TF \xtemp_reg[4]  ( .D(N715), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[8]), .QN(N151) );
  DFFRX2TF \step_reg[3]  ( .D(N721), .CK(CLK), .RN(RST_N), .Q(STEP[3]), .QN(
        N150) );
  DFFRX2TF \step_reg[1]  ( .D(N700), .CK(CLK), .RN(RST_N), .Q(N149), .QN(N121)
         );
  DFFRX2TF \ytemp_reg[12]  ( .D(N706), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[3]), .QN(N148) );
  DFFRX2TF \xtemp_reg[10]  ( .D(N709), .CK(CLK), .RN(RST_N), .Q(XTEMP[10]), 
        .QN(N147) );
  DFFRX2TF \ytemp_reg[8]  ( .D(N686), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_REMA[8]), .QN(N146) );
  DFFRX2TF \xtemp_reg[5]  ( .D(N714), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[9]), .QN(N145) );
  DFFRX2TF \xtemp_reg[3]  ( .D(N716), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[7]), .QN(N144) );
  DFFRX2TF \xtemp_reg[7]  ( .D(N712), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[11]), .QN(N143) );
  DFFRX2TF \step_reg[2]  ( .D(N696), .CK(CLK), .RN(RST_N), .Q(STEP[2]), .QN(
        N142) );
  DFFRX2TF \xtemp_reg[1]  ( .D(N718), .CK(CLK), .RN(RST_N), .Q(
        DIVISION_HEAD[5]), .QN(N141) );
  DFFRX2TF SEL_Z_reg ( .D(N670), .CK(CLK), .RN(RST_N), .Q(N164), .QN(N123) );
  CMPR32X2TF \add_x_132_1/U4  ( .A(OPER_A[10]), .B(OPER_B[10]), .C(
        ADD_X_132_1_N4), .CO(ADD_X_132_1_N3), .S(SUM_AB[10]) );
  CMPR32X2TF \add_x_132_1/U6  ( .A(OPER_A[8]), .B(OPER_B[8]), .C(
        ADD_X_132_1_N6), .CO(ADD_X_132_1_N5), .S(SUM_AB[8]) );
  CMPR32X2TF \add_x_132_1/U8  ( .A(OPER_A[6]), .B(OPER_B[6]), .C(
        ADD_X_132_1_N8), .CO(ADD_X_132_1_N7), .S(SUM_AB[6]) );
  CMPR32X2TF \add_x_132_1/U10  ( .A(OPER_A[4]), .B(OPER_B[4]), .C(
        ADD_X_132_1_N10), .CO(ADD_X_132_1_N9), .S(SUM_AB[4]) );
  CMPR32X2TF \add_x_132_1/U13  ( .A(OPER_A[1]), .B(OPER_B[1]), .C(
        ADD_X_132_1_N13), .CO(ADD_X_132_1_N12), .S(SUM_AB[1]) );
  CMPR32X2TF \add_x_132_1/U5  ( .A(OPER_A[9]), .B(OPER_B[9]), .C(
        ADD_X_132_1_N5), .CO(ADD_X_132_1_N4), .S(SUM_AB[9]) );
  CMPR32X2TF \add_x_132_1/U12  ( .A(OPER_A[2]), .B(OPER_B[2]), .C(
        ADD_X_132_1_N12), .CO(ADD_X_132_1_N11), .S(SUM_AB[2]) );
  CMPR32X2TF \add_x_132_1/U11  ( .A(OPER_A[3]), .B(OPER_B[3]), .C(
        ADD_X_132_1_N11), .CO(ADD_X_132_1_N10), .S(SUM_AB[3]) );
  CMPR32X2TF \add_x_132_1/U9  ( .A(OPER_A[5]), .B(OPER_B[5]), .C(
        ADD_X_132_1_N9), .CO(ADD_X_132_1_N8), .S(SUM_AB[5]) );
  CMPR32X2TF \add_x_132_1/U7  ( .A(OPER_A[7]), .B(OPER_B[7]), .C(
        ADD_X_132_1_N7), .CO(ADD_X_132_1_N6), .S(SUM_AB[7]) );
  CMPR32X2TF \add_x_132_1/U3  ( .A(OPER_A[11]), .B(OPER_B[11]), .C(
        ADD_X_132_1_N3), .CO(ADD_X_132_1_N2), .S(SUM_AB[11]) );
  DFFRX1TF \rsht_bits_reg[2]  ( .D(N701), .CK(CLK), .RN(RST_N), .QN(N90) );
  DFFRX1TF \ztemp_reg[0]  ( .D(N669), .CK(CLK), .RN(RST_N), .Q(ZTEMP[0]) );
  DFFRX1TF \wtemp_reg[6]  ( .D(N676), .CK(CLK), .RN(RST_N), .Q(OPER_B[6]) );
  DFFRX1TF \ztemp_reg[6]  ( .D(N663), .CK(CLK), .RN(RST_N), .Q(ZTEMP[6]) );
  DFFRX1TF \ztemp_reg[4]  ( .D(N665), .CK(CLK), .RN(RST_N), .Q(ZTEMP[4]) );
  DFFRX1TF \ztemp_reg[2]  ( .D(N667), .CK(CLK), .RN(RST_N), .Q(ZTEMP[2]) );
  DFFRX1TF \ztemp_reg[1]  ( .D(N668), .CK(CLK), .RN(RST_N), .Q(ZTEMP[1]) );
  DFFRX1TF \ztemp_reg[5]  ( .D(N664), .CK(CLK), .RN(RST_N), .Q(ZTEMP[5]) );
  DFFRX1TF \ztemp_reg[3]  ( .D(N666), .CK(CLK), .RN(RST_N), .Q(ZTEMP[3]) );
  DFFRX1TF \ztemp_reg[7]  ( .D(N662), .CK(CLK), .RN(RST_N), .Q(ZTEMP[7]) );
  DFFRX1TF \ztemp_reg[8]  ( .D(N661), .CK(CLK), .RN(RST_N), .Q(ZTEMP[8]) );
  DFFRX1TF \ztemp_reg[9]  ( .D(N660), .CK(CLK), .RN(RST_N), .Q(ZTEMP[9]) );
  DFFRX1TF \wtemp_reg[5]  ( .D(N677), .CK(CLK), .RN(RST_N), .Q(OPER_B[5]) );
  DFFRX1TF \wtemp_reg[7]  ( .D(N675), .CK(CLK), .RN(RST_N), .Q(OPER_B[7]) );
  DFFRX1TF \ztemp_reg[10]  ( .D(N659), .CK(CLK), .RN(RST_N), .Q(ZTEMP[10]) );
  DFFRX1TF \ztemp_reg[11]  ( .D(N658), .CK(CLK), .RN(RST_N), .Q(ZTEMP[11]) );
  DFFRX1TF \ztemp_reg[12]  ( .D(N657), .CK(CLK), .RN(RST_N), .Q(ZTEMP[12]) );
  DFFRX2TF XOR_SRC_reg ( .D(N707), .CK(CLK), .RN(RST_N), .Q(N56), .QN(N73) );
  DFFRX2TF \xtemp_reg[9]  ( .D(N710), .CK(CLK), .RN(RST_N), .Q(XTEMP[9]), .QN(
        N529) );
  DFFRX2TF sign_x_reg ( .D(N722), .CK(CLK), .RN(RST_N), .Q(N965), .QN(N74) );
  DFFRX2TF \index_reg[2]  ( .D(N698), .CK(CLK), .RN(RST_N), .Q(\INDEX[2] ) );
  NAND2X1TF U3 ( .A(ALU_START), .B(N259), .Y(N600) );
  AND2X1TF U4 ( .A(N191), .B(ZTEMP[10]), .Y(POUT[10]) );
  OAI222X1TF U5 ( .A0(N87), .A1(N171), .B0(N97), .B1(N147), .C0(N81), .C1(N148), .Y(FOUT[10]) );
  AOI21X1TF U6 ( .A0(N825), .A1(N931), .B0(N848), .Y(N1) );
  NOR3X1TF U7 ( .A(OPER_A[1]), .B(N934), .C(N825), .Y(N2) );
  OAI32X1TF U8 ( .A0(N182), .A1(OPER_B[0]), .A2(N109), .B0(N935), .B1(N182), 
        .Y(N3) );
  AOI211X1TF U9 ( .A0(OPER_B[2]), .A1(N858), .B0(N2), .C0(N3), .Y(N4) );
  OAI31X1TF U10 ( .A0(N109), .A1(N184), .A2(OPER_B[1]), .B0(N824), .Y(N5) );
  AOI211X1TF U11 ( .A0(C152_DATA4_1), .A1(N107), .B0(N886), .C0(N5), .Y(N6) );
  OAI211X1TF U12 ( .A0(N826), .A1(N1), .B0(N4), .C0(N6), .Y(N681) );
  AND2X1TF U13 ( .A(N191), .B(ZTEMP[11]), .Y(POUT[11]) );
  NOR2X1TF U14 ( .A(N98), .B(N155), .Y(FOUT[11]) );
  AOI32X1TF U15 ( .A0(N109), .A1(N837), .A2(N935), .B0(N184), .B1(N837), .Y(N7) );
  AOI211X1TF U16 ( .A0(C152_DATA4_0), .A1(N107), .B0(N886), .C0(N7), .Y(N8) );
  OAI21X1TF U17 ( .A0(N848), .A1(N931), .B0(OPER_A[0]), .Y(N9) );
  OAI211X1TF U18 ( .A0(N182), .A1(N894), .B0(N8), .C0(N9), .Y(N682) );
  NOR3X1TF U19 ( .A(Y_IN[12]), .B(Y_IN[11]), .C(Y_IN[10]), .Y(N10) );
  CLKINVX1TF U20 ( .A(N443), .Y(N11) );
  AOI22X1TF U21 ( .A0(N315), .A1(N11), .B0(N101), .B1(N737), .Y(N12) );
  OAI21X1TF U22 ( .A0(X_IN[4]), .A1(N314), .B0(N85), .Y(N13) );
  OAI22X1TF U23 ( .A0(N101), .A1(N737), .B0(X_IN[6]), .B1(N730), .Y(N14) );
  AOI31X1TF U24 ( .A0(N316), .A1(N12), .A2(N13), .B0(N14), .Y(N15) );
  AOI21X1TF U25 ( .A0(N730), .A1(X_IN[6]), .B0(N15), .Y(N16) );
  OA22X1TF U26 ( .A0(N17), .A1(N16), .B0(N489), .B1(N193), .Y(N18) );
  AO21X1TF U27 ( .A0(N469), .A1(N16), .B0(Y_IN[4]), .Y(N19) );
  AOI22X1TF U28 ( .A0(N489), .A1(N193), .B0(N18), .B1(N19), .Y(N20) );
  AOI2BB2X1TF U29 ( .B0(X_IN[9]), .B1(N20), .A0N(N503), .A1N(N84), .Y(N21) );
  CLKINVX1TF U30 ( .A(N20), .Y(N22) );
  AO21X1TF U31 ( .A0(N501), .A1(N22), .B0(Y_IN[6]), .Y(N23) );
  AOI22X1TF U32 ( .A0(Y_IN[7]), .A1(N503), .B0(N21), .B1(N23), .Y(N24) );
  AOI222XLTF U33 ( .A0(N761), .A1(X_IN[11]), .B0(N761), .B1(N24), .C0(X_IN[11]), .C1(N24), .Y(N25) );
  OAI21X1TF U34 ( .A0(Y_IN[9]), .A1(N302), .B0(N25), .Y(N26) );
  OAI211X1TF U35 ( .A0(X_IN[12]), .A1(N783), .B0(N10), .C0(N26), .Y(N769) );
  CLKINVX1TF U36 ( .A(X_IN[7]), .Y(N17) );
  AND2X1TF U37 ( .A(N191), .B(ZTEMP[12]), .Y(POUT[12]) );
  NOR2X1TF U38 ( .A(N98), .B(N171), .Y(FOUT[12]) );
  AOI22X1TF U39 ( .A0(N117), .A1(ZTEMP[0]), .B0(N1012), .B1(DIVISION_HEAD[0]), 
        .Y(N27) );
  AOI32XLTF U40 ( .A0(N1010), .A1(N27), .A2(N1019), .B0(N976), .B1(N27), .Y(
        N669) );
  OAI32X1TF U41 ( .A0(N185), .A1(N936), .A2(N109), .B0(N935), .B1(N185), .Y(
        N28) );
  CLKINVX1TF U42 ( .A(OPER_A[11]), .Y(N29) );
  OAI32X1TF U43 ( .A0(N29), .A1(N934), .A2(N933), .B0(N932), .B1(N29), .Y(N30)
         );
  AOI31X1TF U44 ( .A0(N933), .A1(N931), .A2(N29), .B0(N930), .Y(N31) );
  NOR2X1TF U45 ( .A(N108), .B(OPER_B[11]), .Y(N32) );
  AOI222XLTF U46 ( .A0(C152_DATA4_11), .A1(N106), .B0(N221), .B1(N964), .C0(
        N936), .C1(N32), .Y(N33) );
  OAI211X1TF U47 ( .A0(N187), .A1(N938), .B0(N31), .C0(N33), .Y(N34) );
  OR3X1TF U48 ( .A(N28), .B(N30), .C(N34), .Y(N671) );
  NOR2X1TF U49 ( .A(N933), .B(OPER_A[11]), .Y(N35) );
  XNOR2X1TF U50 ( .A(OPER_A[12]), .B(N35), .Y(N36) );
  AOI22X1TF U51 ( .A0(N36), .A1(N931), .B0(OPER_A[12]), .B1(N848), .Y(N37) );
  OAI21X1TF U52 ( .A0(N970), .A1(N549), .B0(N133), .Y(N38) );
  XNOR2X1TF U53 ( .A(N38), .B(N78), .Y(N39) );
  XNOR2X1TF U54 ( .A(DP_OP_333_124_4748_N1), .B(N39), .Y(N40) );
  NOR2X1TF U55 ( .A(OPER_B[11]), .B(N936), .Y(N41) );
  OAI31X1TF U56 ( .A0(N108), .A1(N41), .A2(OPER_B[12]), .B0(N824), .Y(N42) );
  AOI211X1TF U57 ( .A0(N107), .A1(N40), .B0(N930), .C0(N42), .Y(N43) );
  OAI31X1TF U58 ( .A0(OPER_B[11]), .A1(N936), .A2(N911), .B0(N868), .Y(N44) );
  AOI32X1TF U59 ( .A0(N120), .A1(OPER_B[12]), .A2(N44), .B0(N218), .B1(
        OPER_B[12]), .Y(N45) );
  NAND4BX1TF U60 ( .AN(N820), .B(N37), .C(N43), .D(N45), .Y(N724) );
  OAI21X1TF U61 ( .A0(N970), .A1(N656), .B0(N202), .Y(N46) );
  CLKMX2X2TF U62 ( .A(N78), .B(DP_OP_333_124_4748_N57), .S0(N46), .Y(
        DP_OP_333_124_4748_N12) );
  XOR2X1TF U63 ( .A(DP_OP_333_124_4748_N57), .B(N46), .Y(C152_DATA4_0) );
  NOR3X1TF U64 ( .A(N910), .B(N74), .C(N907), .Y(N47) );
  NOR2X1TF U65 ( .A(N161), .B(N938), .Y(N48) );
  AOI211X1TF U66 ( .A0(N106), .A1(C152_DATA4_9), .B0(N47), .C0(N48), .Y(N49)
         );
  NOR2X1TF U67 ( .A(N934), .B(OPER_A[9]), .Y(N50) );
  AOI22X1TF U68 ( .A0(SIGN_Y), .A1(N906), .B0(N909), .B1(N50), .Y(N51) );
  OAI21X1TF U69 ( .A0(N109), .A1(N908), .B0(N935), .Y(N52) );
  OAI21X1TF U70 ( .A0(N934), .A1(N909), .B0(N932), .Y(N53) );
  AOI22X1TF U71 ( .A0(OPER_B[9]), .A1(N52), .B0(OPER_A[9]), .B1(N53), .Y(N54)
         );
  NAND3X1TF U72 ( .A(N937), .B(N908), .C(N188), .Y(N55) );
  NAND4X1TF U73 ( .A(N49), .B(N51), .C(N54), .D(N55), .Y(N673) );
  INVX2TF U74 ( .A(N941), .Y(N111) );
  NAND2X2TF U75 ( .A(SIGN_Y), .B(N965), .Y(N971) );
  AOI22X2TF U76 ( .A0(N73), .A1(DIVISION_HEAD[3]), .B0(XTEMP[12]), .B1(N56), 
        .Y(N346) );
  OAI21XLTF U77 ( .A0(N123), .A1(N952), .B0(N951), .Y(N670) );
  NAND2X1TF U78 ( .A(N773), .B(N765), .Y(N396) );
  AND2X2TF U79 ( .A(ZTEMP[4]), .B(N134), .Y(POUT[4]) );
  NOR3BX2TF U80 ( .AN(ALU_TYPE[2]), .B(ALU_TYPE[0]), .C(ALU_TYPE[1]), .Y(N259)
         );
  OA21XLTF U81 ( .A0(SUM_AB[12]), .A1(N650), .B0(N112), .Y(N136) );
  NAND2XLTF U82 ( .A(N799), .B(SUM_AB[8]), .Y(N425) );
  NAND2X1TF U83 ( .A(N929), .B(N203), .Y(N217) );
  AOI2BB1X1TF U84 ( .A0N(N963), .A1N(N962), .B0(N961), .Y(N1011) );
  CLKINVX1TF U85 ( .A(SUM_AB[4]), .Y(N390) );
  AO21X1TF U86 ( .A0(N776), .A1(N373), .B0(N822), .Y(N510) );
  CLKINVX1TF U87 ( .A(N861), .Y(N859) );
  CLKBUFX2TF U88 ( .A(N190), .Y(DP_OP_333_124_4748_N43) );
  AND2XLTF U89 ( .A(\INDEX[2] ), .B(N625), .Y(N311) );
  AND2X2TF U90 ( .A(N191), .B(N73), .Y(N240) );
  AND2X2TF U91 ( .A(N110), .B(N191), .Y(N241) );
  CLKINVX1TF U92 ( .A(N833), .Y(N828) );
  CLKINVX1TF U93 ( .A(N621), .Y(N623) );
  CLKINVX1TF U94 ( .A(N193), .Y(N200) );
  CLKBUFX2TF U95 ( .A(N73), .Y(N972) );
  CLKINVX1TF U96 ( .A(Y_IN[6]), .Y(N199) );
  AOI211X1TF U97 ( .A0(X_IN[3]), .A1(N746), .B0(N441), .C0(N440), .Y(N442) );
  AOI211X1TF U98 ( .A0(X_IN[5]), .A1(N746), .B0(N459), .C0(N458), .Y(N460) );
  AOI211X1TF U99 ( .A0(Y_IN[7]), .A1(N746), .B0(N787), .C0(N786), .Y(N788) );
  OA21XLTF U100 ( .A0(SUM_AB[12]), .A1(N395), .B0(N112), .Y(N506) );
  CLKINVX2TF U101 ( .A(N865), .Y(N211) );
  AOI21X1TF U102 ( .A0(N766), .A1(N306), .B0(N387), .Y(N383) );
  INVX1TF U103 ( .A(N906), .Y(N883) );
  AND2X2TF U104 ( .A(N904), .B(N922), .Y(N937) );
  INVX2TF U105 ( .A(N115), .Y(N116) );
  OAI21XLTF U106 ( .A0(N309), .A1(N629), .B0(N622), .Y(N310) );
  AOI22X1TF U107 ( .A0(X_IN[5]), .A1(N445), .B0(N79), .B1(N99), .Y(N447) );
  OAI31X1TF U108 ( .A0(N282), .A1(X_IN[11]), .A2(N548), .B0(N281), .Y(N283) );
  OAI21X1TF U109 ( .A0(N379), .A1(N746), .B0(N381), .Y(N380) );
  AOI22X1TF U110 ( .A0(Y_IN[9]), .A1(N801), .B0(X_IN[4]), .B1(N131), .Y(N802)
         );
  AOI22X1TF U111 ( .A0(X_IN[2]), .A1(N131), .B0(X_IN[3]), .B1(N806), .Y(N785)
         );
  AOI211X2TF U112 ( .A0(N571), .A1(N941), .B0(N595), .C0(N570), .Y(N597) );
  AOI22X1TF U113 ( .A0(X_IN[12]), .A1(N806), .B0(X_IN[11]), .B1(N131), .Y(N437) );
  INVX1TF U114 ( .A(N405), .Y(N406) );
  AOI21X1TF U115 ( .A0(N643), .A1(N120), .B0(N642), .Y(N646) );
  NAND3XLTF U116 ( .A(N120), .B(N823), .C(N822), .Y(N633) );
  OAI31X1TF U117 ( .A0(N565), .A1(N566), .A2(N564), .B0(N120), .Y(N582) );
  AOI22X1TF U118 ( .A0(XTEMP[11]), .A1(N126), .B0(N79), .B1(N445), .Y(N354) );
  AOI32XLTF U119 ( .A0(N821), .A1(N941), .A2(N822), .B0(N638), .B1(N120), .Y(
        N644) );
  OAI2BB2XLTF U120 ( .B0(N761), .B1(N803), .A0N(Y_IN[6]), .A1N(N801), .Y(N778)
         );
  OAI31XLTF U121 ( .A0(N112), .A1(N165), .A2(N632), .B0(N631), .Y(N637) );
  OR2X2TF U122 ( .A(N387), .B(N763), .Y(N800) );
  NAND4XLTF U123 ( .A(N612), .B(N611), .C(N610), .D(N609), .Y(N613) );
  AOI22X1TF U124 ( .A0(Y_IN[1]), .A1(N801), .B0(DIVISION_REMA[4]), .B1(N114), 
        .Y(N731) );
  INVX1TF U125 ( .A(OPER_A[1]), .Y(N826) );
  INVX1TF U126 ( .A(OPER_A[0]), .Y(N825) );
  AOI22X1TF U127 ( .A0(XTEMP[10]), .A1(N88), .B0(X_IN[7]), .B1(N801), .Y(N481)
         );
  INVX1TF U128 ( .A(OPER_A[10]), .Y(N915) );
  AOI22X1TF U129 ( .A0(DIVISION_HEAD[2]), .A1(N114), .B0(Y_IN[8]), .B1(N801), 
        .Y(N794) );
  OAI211XLTF U130 ( .A0(N970), .A1(N365), .B0(N973), .C0(N601), .Y(N367) );
  NAND3BXLTF U131 ( .AN(N382), .B(N776), .C(N639), .Y(N366) );
  INVX1TF U132 ( .A(OPER_A[8]), .Y(N897) );
  AOI22X1TF U133 ( .A0(N193), .A1(N801), .B0(Y_IN[7]), .B1(N790), .Y(N754) );
  INVX1TF U134 ( .A(OPER_A[4]), .Y(N856) );
  AOI22X1TF U135 ( .A0(Y_IN[3]), .A1(N801), .B0(DIVISION_REMA[6]), .B1(N114), 
        .Y(N741) );
  AOI22X1TF U136 ( .A0(X_IN[2]), .A1(N801), .B0(X_IN[3]), .B1(N445), .Y(N426)
         );
  INVX1TF U137 ( .A(OPER_A[6]), .Y(N875) );
  AOI22X1TF U138 ( .A0(DIVISION_HEAD[3]), .A1(N103), .B0(ZTEMP[12]), .B1(N135), 
        .Y(N256) );
  AOI22X1TF U139 ( .A0(DIVISION_REMA[8]), .A1(N103), .B0(ZTEMP[8]), .B1(N164), 
        .Y(N251) );
  INVX2TF U140 ( .A(N735), .Y(N93) );
  AOI22X1TF U141 ( .A0(DIVISION_HEAD[2]), .A1(N103), .B0(ZTEMP[11]), .B1(N135), 
        .Y(N254) );
  AOI22X1TF U142 ( .A0(DIVISION_HEAD[0]), .A1(N103), .B0(ZTEMP[9]), .B1(N135), 
        .Y(N252) );
  AOI22X1TF U143 ( .A0(DIVISION_REMA[7]), .A1(N103), .B0(ZTEMP[7]), .B1(N164), 
        .Y(N250) );
  AOI22X1TF U144 ( .A0(DIVISION_HEAD[1]), .A1(N103), .B0(ZTEMP[10]), .B1(N135), 
        .Y(N253) );
  AOI22X1TF U145 ( .A0(DIVISION_REMA[5]), .A1(N103), .B0(ZTEMP[5]), .B1(N164), 
        .Y(N248) );
  AOI22X1TF U146 ( .A0(DIVISION_REMA[6]), .A1(N103), .B0(ZTEMP[6]), .B1(N164), 
        .Y(N249) );
  INVX2TF U147 ( .A(DP_OP_333_124_4748_N43), .Y(N78) );
  INVX2TF U148 ( .A(N746), .Y(N95) );
  AOI22X1TF U149 ( .A0(DIVISION_REMA[4]), .A1(N103), .B0(ZTEMP[4]), .B1(N164), 
        .Y(N247) );
  AOI22X1TF U150 ( .A0(DIVISION_REMA[3]), .A1(N103), .B0(ZTEMP[3]), .B1(N164), 
        .Y(N246) );
  AOI22X1TF U151 ( .A0(DIVISION_REMA[0]), .A1(N102), .B0(ZTEMP[0]), .B1(N164), 
        .Y(N243) );
  AOI22X1TF U152 ( .A0(DIVISION_REMA[2]), .A1(N102), .B0(ZTEMP[2]), .B1(N164), 
        .Y(N245) );
  AOI22X1TF U153 ( .A0(DIVISION_REMA[1]), .A1(N102), .B0(ZTEMP[1]), .B1(N164), 
        .Y(N244) );
  INVX2TF U154 ( .A(N255), .Y(N102) );
  OAI21XLTF U155 ( .A0(N970), .A1(N314), .B0(N202), .Y(C2_Z_1) );
  CLKAND2X2TF U156 ( .A(N647), .B(N640), .Y(N546) );
  INVX2TF U157 ( .A(N812), .Y(N113) );
  NAND2BXLTF U158 ( .AN(DP_OP_333_124_4748_N57), .B(N970), .Y(N203) );
  AND2X2TF U159 ( .A(N384), .B(N351), .Y(N735) );
  AND2X2TF U160 ( .A(N342), .B(N219), .Y(N941) );
  AND2X2TF U161 ( .A(N351), .B(DP_OP_333_124_4748_N57), .Y(N746) );
  INVX1TF U162 ( .A(N342), .Y(N955) );
  NAND2XLTF U163 ( .A(N219), .B(N946), .Y(N534) );
  AND2X2TF U164 ( .A(N123), .B(N242), .Y(N257) );
  OR2X2TF U165 ( .A(N164), .B(N242), .Y(N255) );
  OR3X1TF U166 ( .A(PRE_WORK), .B(N606), .C(N600), .Y(N502) );
  OR2X2TF U167 ( .A(N348), .B(N600), .Y(N812) );
  CLKAND2X2TF U168 ( .A(ZTEMP[2]), .B(N134), .Y(POUT[2]) );
  CLKAND2X2TF U169 ( .A(ZTEMP[5]), .B(N134), .Y(POUT[5]) );
  CLKAND2X2TF U170 ( .A(ZTEMP[3]), .B(N134), .Y(POUT[3]) );
  CLKAND2X2TF U171 ( .A(ZTEMP[9]), .B(N134), .Y(POUT[9]) );
  CLKAND2X2TF U172 ( .A(ZTEMP[1]), .B(N134), .Y(POUT[1]) );
  INVX2TF U173 ( .A(N972), .Y(N110) );
  INVX2TF U174 ( .A(N196), .Y(N101) );
  CLKAND2X2TF U175 ( .A(ZTEMP[7]), .B(N191), .Y(POUT[7]) );
  CLKAND2X2TF U176 ( .A(ZTEMP[6]), .B(N191), .Y(POUT[6]) );
  CLKAND2X2TF U177 ( .A(ZTEMP[0]), .B(N191), .Y(POUT[0]) );
  INVX2TF U178 ( .A(N194), .Y(N84) );
  CLKAND2X2TF U179 ( .A(ZTEMP[8]), .B(N191), .Y(POUT[8]) );
  NAND2XLTF U180 ( .A(DIVISION_HEAD[4]), .B(N259), .Y(N222) );
  AOI22X1TF U181 ( .A0(X_IN[11]), .A1(N548), .B0(X_IN[12]), .B1(N804), .Y(N277) );
  INVX2TF U182 ( .A(X_IN[3]), .Y(N195) );
  INVX2TF U183 ( .A(X_IN[5]), .Y(N196) );
  INVX1TF U184 ( .A(X_IN[2]), .Y(N771) );
  INVX2TF U185 ( .A(Y_IN[7]), .Y(N194) );
  INVX2TF U186 ( .A(N298), .Y(N79) );
  INVX2TF U187 ( .A(N241), .Y(N80) );
  INVX2TF U188 ( .A(N241), .Y(N81) );
  INVX2TF U189 ( .A(N1019), .Y(N82) );
  INVX2TF U190 ( .A(N1019), .Y(N83) );
  INVX2TF U191 ( .A(N195), .Y(N85) );
  INVX2TF U192 ( .A(N240), .Y(N86) );
  INVX2TF U193 ( .A(N240), .Y(N87) );
  INVX2TF U194 ( .A(N502), .Y(N88) );
  INVX2TF U195 ( .A(N502), .Y(N89) );
  INVX2TF U196 ( .A(N735), .Y(N94) );
  INVX2TF U197 ( .A(N746), .Y(N96) );
  INVX2TF U198 ( .A(N259), .Y(N97) );
  INVX2TF U199 ( .A(N259), .Y(N98) );
  INVX2TF U200 ( .A(N396), .Y(N99) );
  INVX2TF U201 ( .A(N396), .Y(N100) );
  INVX2TF U202 ( .A(N255), .Y(N103) );
  INVX2TF U203 ( .A(N257), .Y(N104) );
  INVX2TF U204 ( .A(N257), .Y(N105) );
  INVX2TF U205 ( .A(N217), .Y(N106) );
  INVX2TF U206 ( .A(N217), .Y(N107) );
  INVX2TF U207 ( .A(N937), .Y(N108) );
  INVX2TF U208 ( .A(N937), .Y(N109) );
  INVX2TF U209 ( .A(N941), .Y(N112) );
  INVX2TF U210 ( .A(N812), .Y(N114) );
  INVX2TF U211 ( .A(N1011), .Y(N115) );
  INVX2TF U212 ( .A(N115), .Y(N117) );
  INVX2TF U213 ( .A(N510), .Y(N118) );
  INVX2TF U214 ( .A(N510), .Y(N119) );
  INVX2TF U215 ( .A(N111), .Y(N120) );
  INVX2TF U216 ( .A(DP_OP_333_124_4748_N43), .Y(N125) );
  INVX2TF U217 ( .A(N93), .Y(N126) );
  AOI222X4TF U218 ( .A0(N488), .A1(N147), .B0(N488), .B1(N503), .C0(N147), 
        .C1(N503), .Y(N498) );
  NOR2X2TF U219 ( .A(N339), .B(N956), .Y(N351) );
  NOR2X2TF U220 ( .A(N348), .B(N970), .Y(N384) );
  NOR3X2TF U221 ( .A(N111), .B(N605), .C(N632), .Y(N618) );
  INVX2TF U222 ( .A(N506), .Y(N127) );
  INVX2TF U223 ( .A(N506), .Y(N130) );
  INVX2TF U224 ( .A(N800), .Y(N131) );
  INVX2TF U225 ( .A(N800), .Y(N132) );
  NAND2X2TF U226 ( .A(N123), .B(N762), .Y(N455) );
  AOI21X2TF U227 ( .A0(N941), .A1(N921), .B0(N218), .Y(N935) );
  AOI211XLTF U228 ( .A0(N826), .A1(N825), .B0(OPER_A[2]), .C0(N916), .Y(N827)
         );
  OAI32XLTF U229 ( .A0(OPER_A[8]), .A1(N898), .A2(N916), .B0(N897), .B1(N896), 
        .Y(N899) );
  OAI32XLTF U230 ( .A0(OPER_A[10]), .A1(N917), .A2(N916), .B0(N915), .B1(N914), 
        .Y(N918) );
  OAI32XLTF U231 ( .A0(OPER_A[6]), .A1(N876), .A2(N916), .B0(N875), .B1(N874), 
        .Y(N877) );
  INVXLTF U232 ( .A(N916), .Y(N913) );
  INVX2TF U233 ( .A(DP_OP_333_124_4748_N57), .Y(N133) );
  CLKBUFX2TF U234 ( .A(N191), .Y(N134) );
  CLKBUFX2TF U235 ( .A(N258), .Y(N191) );
  NOR3XLTF U236 ( .A(N73), .B(N910), .C(N971), .Y(N820) );
  NAND2X2TF U237 ( .A(N969), .B(N929), .Y(N910) );
  AOI21XLTF U238 ( .A0(N821), .A1(N375), .B0(N374), .Y(N377) );
  AOI21XLTF U239 ( .A0(N823), .A1(N822), .B0(N821), .Y(N829) );
  INVXLTF U240 ( .A(N821), .Y(N378) );
  NOR3BX4TF U241 ( .AN(N386), .B(N383), .C(N126), .Y(N514) );
  AOI222X4TF U242 ( .A0(XTEMP[9]), .A1(X_IN[9]), .B0(XTEMP[9]), .B1(N479), 
        .C0(X_IN[9]), .C1(N479), .Y(N488) );
  AOI222X4TF U243 ( .A0(N176), .A1(N489), .B0(N176), .B1(N465), .C0(N489), 
        .C1(N465), .Y(N479) );
  OAI31XLTF U244 ( .A0(OPER_A[1]), .A1(N916), .A2(OPER_A[0]), .B0(N831), .Y(
        N832) );
  OAI21X2TF U245 ( .A0(N141), .A1(N104), .B0(N244), .Y(OPER_A[1]) );
  INVX2TF U246 ( .A(N123), .Y(N135) );
  NAND2X2TF U247 ( .A(N762), .B(N135), .Y(N559) );
  NOR2X4TF U248 ( .A(N387), .B(N768), .Y(N806) );
  AOI22XLTF U249 ( .A0(DIVISION_HEAD[5]), .A1(N88), .B0(X_IN[7]), .B1(N806), 
        .Y(N389) );
  AOI22XLTF U250 ( .A0(X_IN[10]), .A1(N131), .B0(X_IN[11]), .B1(N806), .Y(N428) );
  NOR4X2TF U251 ( .A(N648), .B(N943), .C(N367), .D(N366), .Y(N642) );
  NOR2X2TF U252 ( .A(N339), .B(N604), .Y(N566) );
  NOR2BX2TF U253 ( .AN(N544), .B(N384), .Y(N629) );
  INVX2TF U254 ( .A(N136), .Y(N137) );
  INVX2TF U255 ( .A(N136), .Y(N138) );
  AOI22X2TF U256 ( .A0(N346), .A1(N344), .B0(N940), .B1(N347), .Y(N922) );
  CLKBUFX2TF U257 ( .A(N1012), .Y(N139) );
  NOR2X1TF U258 ( .A(N116), .B(N190), .Y(N1012) );
  XNOR2X1TF U259 ( .A(OPER_A[12]), .B(ADD_X_132_1_N2), .Y(N140) );
  XNOR2X2TF U260 ( .A(N140), .B(OPER_B[12]), .Y(SUM_AB[12]) );
  ADDHX1TF U261 ( .A(OPER_B[0]), .B(OPER_A[0]), .CO(ADD_X_132_1_N13), .S(
        SUM_AB[0]) );
  AOI222XLTF U262 ( .A0(DIVISION_HEAD[1]), .A1(DIVISION_HEAD[0]), .B0(
        DIVISION_HEAD[1]), .B1(N315), .C0(DIVISION_HEAD[0]), .C1(N314), .Y(
        N317) );
  NAND2X1TF U263 ( .A(N314), .B(N656), .Y(N316) );
  AOI22X1TF U264 ( .A0(N73), .A1(N162), .B0(POST_WORK), .B1(N110), .Y(N242) );
  OAI31X1TF U265 ( .A0(N970), .A1(N949), .A2(N948), .B0(N947), .Y(N950) );
  INVX2TF U266 ( .A(N929), .Y(N218) );
  OAI21X1TF U267 ( .A0(N948), .A1(N610), .B0(N647), .Y(N961) );
  NAND2X1TF U268 ( .A(N478), .B(N477), .Y(N487) );
  NOR2X1TF U269 ( .A(SUM_AB[8]), .B(N463), .Y(N478) );
  OA22X1TF U270 ( .A0(N768), .A1(N558), .B0(N763), .B1(N764), .Y(N306) );
  NAND2X1TF U271 ( .A(Y_IN[1]), .B(Y_IN[0]), .Y(N315) );
  NAND2X1TF U272 ( .A(N565), .B(N347), .Y(N916) );
  NOR2X2TF U273 ( .A(N218), .B(N111), .Y(N904) );
  OR2X2TF U274 ( .A(N961), .B(N198), .Y(N929) );
  OAI21X1TF U275 ( .A0(DIVISION_HEAD[12]), .A1(N549), .B0(N338), .Y(N948) );
  AOI2BB1X1TF U276 ( .A0N(DIVISION_HEAD[6]), .A1N(N327), .B0(Y_IN[6]), .Y(N325) );
  AOI2BB1X1TF U277 ( .A0N(DIVISION_HEAD[4]), .A1N(N323), .B0(Y_IN[4]), .Y(N321) );
  NOR2X1TF U278 ( .A(SUM_AB[10]), .B(N487), .Y(N500) );
  NOR2X1TF U279 ( .A(\INDEX[2] ), .B(N621), .Y(N309) );
  NAND2X1TF U280 ( .A(N129), .B(N128), .Y(N621) );
  NAND2X1TF U281 ( .A(N912), .B(N904), .Y(N932) );
  AOI2BB1X1TF U282 ( .A0N(N608), .A1N(N343), .B0(N962), .Y(N198) );
  NAND2X1TF U283 ( .A(PRE_WORK), .B(N125), .Y(N387) );
  CLKBUFX2TF U284 ( .A(N970), .Y(N190) );
  AOI211X1TF U285 ( .A0(Y_IN[11]), .A1(N302), .B0(Y_IN[12]), .C0(N283), .Y(
        N766) );
  CLKBUFX2TF U286 ( .A(Y_IN[5]), .Y(N193) );
  NOR2X1TF U287 ( .A(PRE_WORK), .B(N340), .Y(N342) );
  NOR2X1TF U288 ( .A(N124), .B(N628), .Y(N340) );
  NAND2X1TF U289 ( .A(N122), .B(N149), .Y(N605) );
  NAND2X1TF U290 ( .A(N175), .B(N365), .Y(N348) );
  NAND2X1TF U291 ( .A(N142), .B(N150), .Y(N339) );
  NAND2X1TF U292 ( .A(N455), .B(N461), .Y(N472) );
  NAND2X2TF U293 ( .A(N547), .B(N386), .Y(N461) );
  NAND2X1TF U294 ( .A(N566), .B(N384), .Y(N610) );
  NAND2X1TF U295 ( .A(N121), .B(N165), .Y(N604) );
  CLKBUFX2TF U296 ( .A(N781), .Y(N192) );
  NAND2X1TF U297 ( .A(N121), .B(N122), .Y(N956) );
  AND2X2TF U298 ( .A(ALU_START), .B(N134), .Y(N219) );
  NAND2X2TF U299 ( .A(N220), .B(ALU_START), .Y(N970) );
  NAND2X1TF U300 ( .A(N124), .B(N309), .Y(N365) );
  AND2X2TF U301 ( .A(N197), .B(ALU_TYPE[1]), .Y(N220) );
  AOI211X1TF U302 ( .A0(N219), .A1(N608), .B0(N945), .C0(N607), .Y(N611) );
  NOR3X1TF U303 ( .A(N606), .B(N605), .C(N776), .Y(N607) );
  OR3X1TF U304 ( .A(N882), .B(N881), .C(N213), .Y(N676) );
  OAI2BB2XLTF U305 ( .B0(N883), .B1(N971), .A0N(C152_DATA4_6), .A1N(N107), .Y(
        N213) );
  OAI2BB2XLTF U306 ( .B0(N880), .B1(N924), .A0N(N218), .A1N(OPER_B[6]), .Y(
        N881) );
  AOI32X1TF U307 ( .A0(N969), .A1(N115), .A2(N968), .B0(N120), .B1(N115), .Y(
        N1019) );
  INVX2TF U308 ( .A(N461), .Y(N476) );
  NAND2X1TF U309 ( .A(N904), .B(N871), .Y(N894) );
  NOR2X1TF U310 ( .A(N56), .B(N910), .Y(N906) );
  AOI21X1TF U311 ( .A0(N949), .A1(N967), .B0(N363), .Y(N969) );
  NAND2X1TF U312 ( .A(N340), .B(N175), .Y(N345) );
  NOR2BX2TF U313 ( .AN(N547), .B(N557), .Y(N813) );
  NAND2X1TF U314 ( .A(N142), .B(STEP[3]), .Y(N632) );
  NOR2X1TF U315 ( .A(N175), .B(N600), .Y(N353) );
  NAND3X1TF U316 ( .A(N962), .B(N970), .C(N600), .Y(N647) );
  INVX2TF U317 ( .A(N219), .Y(N962) );
  NAND2X1TF U318 ( .A(N960), .B(DP_OP_333_124_4748_N57), .Y(N650) );
  AND2X2TF U319 ( .A(N219), .B(PRE_WORK), .Y(DP_OP_333_124_4748_N57) );
  INVX2TF U320 ( .A(N364), .Y(N762) );
  NAND2X1TF U321 ( .A(N384), .B(N960), .Y(N364) );
  NOR2X2TF U322 ( .A(N339), .B(N605), .Y(N960) );
  NOR3BX1TF U323 ( .AN(ALU_TYPE[0]), .B(ALU_TYPE[1]), .C(ALU_TYPE[2]), .Y(N258) );
  AO22X1TF U324 ( .A0(N372), .A1(XTEMP[12]), .B0(N360), .B1(N965), .Y(N722) );
  AOI32X1TF U325 ( .A0(N967), .A1(N361), .A2(N958), .B0(N973), .B1(N361), .Y(
        N362) );
  NAND2X1TF U326 ( .A(N946), .B(DP_OP_333_124_4748_N57), .Y(N635) );
  NAND2X1TF U327 ( .A(N643), .B(N114), .Y(N615) );
  NAND2X1TF U328 ( .A(N107), .B(C152_DATA4_8), .Y(N214) );
  AOI32X1TF U329 ( .A0(N118), .A1(DIVISION_HEAD[4]), .A2(N749), .B0(N472), 
        .B1(DIVISION_HEAD[4]), .Y(N393) );
  OAI22X1TF U330 ( .A0(N529), .A1(N94), .B0(N489), .B1(N96), .Y(N490) );
  INVX2TF U331 ( .A(N1015), .Y(N1010) );
  OAI2BB2XLTF U332 ( .B0(N56), .B1(N971), .A0N(N971), .A1N(N56), .Y(N974) );
  NAND2X1TF U333 ( .A(N647), .B(N95), .Y(N944) );
  NAND2X1TF U334 ( .A(N566), .B(DP_OP_333_124_4748_N57), .Y(N395) );
  NOR2X1TF U335 ( .A(N605), .B(N954), .Y(N565) );
  NAND2X1TF U336 ( .A(STEP[2]), .B(N150), .Y(N954) );
  INVX2TF U337 ( .A(N113), .Y(N776) );
  NOR2X2TF U338 ( .A(N762), .B(N192), .Y(N760) );
  NAND2X1TF U339 ( .A(N351), .B(N113), .Y(N544) );
  NOR2X1TF U340 ( .A(N956), .B(N632), .Y(N564) );
  OAI21X2TF U341 ( .A0(N153), .A1(N104), .B0(N243), .Y(OPER_A[0]) );
  OAI32X1TF U342 ( .A0(N649), .A1(N178), .A2(N944), .B0(N148), .B1(N650), .Y(
        N694) );
  OAI21X1TF U343 ( .A0(N175), .A1(N648), .B0(N647), .Y(N695) );
  AOI22X1TF U344 ( .A0(N543), .A1(N73), .B0(N542), .B1(N541), .Y(N707) );
  INVX2TF U345 ( .A(N543), .Y(N541) );
  OAI31X1TF U346 ( .A0(N540), .A1(N539), .A2(N538), .B0(N537), .Y(N542) );
  AOI211X1TF U347 ( .A0(N536), .A1(XTEMP[12]), .B0(N535), .C0(N534), .Y(N537)
         );
  OAI31X1TF U348 ( .A0(DIVISION_HEAD[1]), .A1(N533), .A2(N147), .B0(N532), .Y(
        N536) );
  AOI22X1TF U349 ( .A0(N531), .A1(N530), .B0(XTEMP[11]), .B1(N163), .Y(N532)
         );
  OAI22X1TF U350 ( .A0(DIVISION_HEAD[0]), .A1(N529), .B0(DIVISION_REMA[8]), 
        .B1(N176), .Y(N530) );
  INVX2TF U351 ( .A(N539), .Y(N531) );
  NOR2X1TF U352 ( .A(XTEMP[11]), .B(N163), .Y(N533) );
  OAI22X1TF U353 ( .A0(DIVISION_HEAD[12]), .A1(N146), .B0(XTEMP[12]), .B1(N148), .Y(N538) );
  OAI21X1TF U354 ( .A0(XTEMP[11]), .A1(N163), .B0(N528), .Y(N539) );
  AOI22X1TF U355 ( .A0(DIVISION_HEAD[0]), .A1(N529), .B0(DIVISION_HEAD[1]), 
        .B1(N147), .Y(N528) );
  AOI21X1TF U356 ( .A0(DIVISION_HEAD[11]), .A1(N168), .B0(N527), .Y(N540) );
  AOI211X1TF U357 ( .A0(DIVISION_REMA[6]), .A1(N154), .B0(N526), .C0(N525), 
        .Y(N527) );
  NOR2X1TF U358 ( .A(DIVISION_HEAD[11]), .B(N168), .Y(N525) );
  AOI21X1TF U359 ( .A0(DIVISION_HEAD[9]), .A1(N167), .B0(N523), .Y(N524) );
  AOI211X1TF U360 ( .A0(DIVISION_REMA[4]), .A1(N151), .B0(N522), .C0(N521), 
        .Y(N523) );
  NOR2X1TF U361 ( .A(DIVISION_HEAD[9]), .B(N167), .Y(N521) );
  AOI21X1TF U362 ( .A0(DIVISION_HEAD[7]), .A1(N166), .B0(N519), .Y(N520) );
  AOI211X1TF U363 ( .A0(N518), .A1(DIVISION_REMA[2]), .B0(N517), .C0(N516), 
        .Y(N519) );
  NOR2X1TF U364 ( .A(DIVISION_HEAD[7]), .B(N166), .Y(N517) );
  OAI21X1TF U365 ( .A0(DIVISION_HEAD[5]), .A1(N159), .B0(N515), .Y(N518) );
  OAI211X1TF U366 ( .A0(DIVISION_REMA[1]), .A1(N141), .B0(DIVISION_REMA[0]), 
        .C0(N153), .Y(N515) );
  OAI21X1TF U367 ( .A0(N381), .A1(N162), .B0(N380), .Y(N720) );
  OAI22X1TF U368 ( .A0(N112), .A1(N378), .B0(N763), .B1(N640), .Y(N379) );
  OAI211X1TF U369 ( .A0(N373), .A1(N822), .B0(N612), .C0(N640), .Y(N374) );
  OAI21X1TF U370 ( .A0(N950), .A1(N969), .B0(N952), .Y(N951) );
  OR4X2TF U371 ( .A(N945), .B(N944), .C(N943), .D(N942), .Y(N952) );
  OAI22X1TF U372 ( .A0(N112), .A1(N940), .B0(N939), .B1(N973), .Y(N942) );
  OAI21X1TF U373 ( .A0(N597), .A1(N586), .B0(N585), .Y(N702) );
  AOI31X1TF U374 ( .A0(N584), .A1(N589), .A2(N591), .B0(N583), .Y(N586) );
  OAI22X1TF U375 ( .A0(N128), .A1(N582), .B0(N593), .B1(N589), .Y(N583) );
  OAI21X1TF U376 ( .A0(N128), .A1(N620), .B0(N619), .Y(N699) );
  AOI31X1TF U377 ( .A0(N618), .A1(N621), .A2(N617), .B0(N616), .Y(N619) );
  OAI32X1TF U378 ( .A0(N629), .A1(N630), .A2(N621), .B0(N617), .B1(N629), .Y(
        N616) );
  AOI22X1TF U379 ( .A0(N597), .A1(N92), .B0(N581), .B1(N580), .Y(N703) );
  AOI211X1TF U380 ( .A0(N595), .A1(N157), .B0(N579), .C0(N790), .Y(N581) );
  AOI21X1TF U381 ( .A0(N578), .A1(N776), .B0(N180), .Y(N579) );
  OAI21X1TF U382 ( .A0(N129), .A1(N620), .B0(N308), .Y(N726) );
  OAI21X1TF U383 ( .A0(N307), .A1(N383), .B0(N620), .Y(N308) );
  AOI32X1TF U384 ( .A0(N629), .A1(N635), .A2(N376), .B0(N157), .B1(N635), .Y(
        N307) );
  OAI31X1TF U385 ( .A0(N630), .A1(N629), .A2(N628), .B0(N627), .Y(N698) );
  AOI22X1TF U386 ( .A0(\INDEX[2] ), .A1(N626), .B0(N625), .B1(N624), .Y(N627)
         );
  OAI21X1TF U387 ( .A0(N623), .A1(N629), .B0(N622), .Y(N626) );
  AOI32X1TF U388 ( .A0(N311), .A1(N124), .A2(N618), .B0(N186), .B1(N310), .Y(
        N313) );
  NOR2X1TF U389 ( .A(N630), .B(N624), .Y(N622) );
  AOI21X1TF U390 ( .A0(\INDEX[2] ), .A1(N625), .B0(N376), .Y(N624) );
  INVX2TF U391 ( .A(N620), .Y(N630) );
  INVX2TF U392 ( .A(N617), .Y(N625) );
  OAI211X1TF U393 ( .A0(N112), .A1(N369), .B0(N645), .C0(N368), .Y(N721) );
  AOI22X1TF U394 ( .A0(STEP[3]), .A1(N642), .B0(N375), .B1(N574), .Y(N368) );
  OAI211X1TF U395 ( .A0(N179), .A1(N615), .B0(N631), .C0(N614), .Y(N700) );
  AOI21X1TF U396 ( .A0(N642), .A1(N149), .B0(N613), .Y(N614) );
  NOR3X1TF U397 ( .A(STEP[3]), .B(N112), .C(N604), .Y(N945) );
  AOI211X1TF U398 ( .A0(N823), .A1(N375), .B0(N372), .C0(N371), .Y(N612) );
  AOI21X1TF U399 ( .A0(N385), .A1(N370), .B0(N776), .Y(N371) );
  NOR2X1TF U400 ( .A(N111), .B(N822), .Y(N375) );
  OAI22X1TF U401 ( .A0(N90), .A1(N598), .B0(N597), .B1(N596), .Y(N701) );
  AOI21X1TF U402 ( .A0(\INDEX[2] ), .A1(N595), .B0(N594), .Y(N596) );
  OAI22X1TF U403 ( .A0(N593), .A1(N592), .B0(N591), .B1(N590), .Y(N594) );
  INVX2TF U404 ( .A(N588), .Y(N593) );
  AOI21X1TF U405 ( .A0(N589), .A1(N588), .B0(N587), .Y(N598) );
  OAI211X1TF U406 ( .A0(N646), .A1(N142), .B0(N645), .C0(N644), .Y(N696) );
  NOR2X1TF U407 ( .A(N649), .B(N362), .Y(N645) );
  OAI21X1TF U408 ( .A0(N351), .A1(N260), .B0(N120), .Y(N361) );
  INVX2TF U409 ( .A(N650), .Y(N649) );
  OAI22X1TF U410 ( .A0(N165), .A1(N954), .B0(N822), .B1(N967), .Y(N638) );
  AOI211X1TF U411 ( .A0(N642), .A1(N165), .B0(N637), .C0(N636), .Y(N641) );
  INVX2TF U412 ( .A(N261), .Y(N634) );
  AOI31X1TF U413 ( .A0(N956), .A1(N370), .A2(N385), .B0(N776), .Y(N261) );
  AOI21X1TF U414 ( .A0(N125), .A1(N603), .B0(N602), .Y(N631) );
  OAI21X1TF U415 ( .A0(N601), .A1(N600), .B0(N599), .Y(N602) );
  OAI22X1TF U416 ( .A0(N597), .A1(N577), .B0(N576), .B1(N189), .Y(N704) );
  AOI21X1TF U417 ( .A0(N592), .A1(N588), .B0(N587), .Y(N576) );
  OAI21X1TF U418 ( .A0(N90), .A1(N591), .B0(N584), .Y(N590) );
  INVX2TF U419 ( .A(N615), .Y(N584) );
  INVX2TF U420 ( .A(N597), .Y(N580) );
  OAI31X1TF U421 ( .A0(N606), .A1(N605), .A2(N776), .B0(N578), .Y(N588) );
  OAI32X1TF U422 ( .A0(N575), .A1(N823), .A2(N574), .B0(N120), .B1(N575), .Y(
        N578) );
  INVX2TF U423 ( .A(N573), .Y(N575) );
  AOI21X1TF U424 ( .A0(N595), .A1(N186), .B0(N572), .Y(N577) );
  AOI32X1TF U425 ( .A0(N566), .A1(N114), .A2(N179), .B0(N960), .B1(N113), .Y(
        N568) );
  AOI31X1TF U426 ( .A0(N120), .A1(N823), .A2(N822), .B0(N944), .Y(N569) );
  INVX2TF U427 ( .A(N582), .Y(N595) );
  AOI22X1TF U428 ( .A0(N903), .A1(N904), .B0(N218), .B1(OPER_B[8]), .Y(N215)
         );
  OAI21X1TF U429 ( .A0(N902), .A1(N160), .B0(N901), .Y(N903) );
  AOI211X1TF U430 ( .A0(N920), .A1(OPER_B[9]), .B0(N900), .C0(N899), .Y(N901)
         );
  AOI21X1TF U431 ( .A0(N913), .A1(N898), .B0(N912), .Y(N896) );
  NOR3X1TF U432 ( .A(N911), .B(OPER_B[8]), .C(N895), .Y(N900) );
  AOI21X1TF U433 ( .A0(N895), .A1(N922), .B0(N921), .Y(N902) );
  OAI211X1TF U434 ( .A0(N1010), .A1(N991), .B0(N990), .C0(N989), .Y(N664) );
  AOI22X1TF U435 ( .A0(DIVISION_HEAD[5]), .A1(N139), .B0(ZTEMP[5]), .B1(N117), 
        .Y(N990) );
  OAI211X1TF U436 ( .A0(N1010), .A1(N997), .B0(N996), .C0(N995), .Y(N662) );
  AOI22X1TF U437 ( .A0(DIVISION_HEAD[7]), .A1(N1012), .B0(ZTEMP[7]), .B1(N117), 
        .Y(N996) );
  OAI211X1TF U438 ( .A0(N1010), .A1(N985), .B0(N984), .C0(N983), .Y(N666) );
  AOI22X1TF U439 ( .A0(DIVISION_HEAD[3]), .A1(N139), .B0(ZTEMP[3]), .B1(N117), 
        .Y(N984) );
  AOI22X1TF U440 ( .A0(SUM_AB[6]), .A1(N82), .B0(N992), .B1(N1015), .Y(N993)
         );
  AOI22X1TF U441 ( .A0(DIVISION_HEAD[6]), .A1(N139), .B0(ZTEMP[6]), .B1(N117), 
        .Y(N994) );
  AOI22X1TF U442 ( .A0(SUM_AB[2]), .A1(N82), .B0(N980), .B1(N1015), .Y(N981)
         );
  AOI22X1TF U443 ( .A0(DIVISION_HEAD[2]), .A1(N139), .B0(ZTEMP[2]), .B1(N116), 
        .Y(N982) );
  AOI22X1TF U444 ( .A0(SUM_AB[4]), .A1(N82), .B0(N986), .B1(N1015), .Y(N987)
         );
  AOI22X1TF U445 ( .A0(DIVISION_HEAD[4]), .A1(N139), .B0(ZTEMP[4]), .B1(N116), 
        .Y(N988) );
  AOI22X1TF U446 ( .A0(SUM_AB[1]), .A1(N82), .B0(N977), .B1(N1015), .Y(N978)
         );
  AOI22X1TF U447 ( .A0(DIVISION_HEAD[1]), .A1(N139), .B0(ZTEMP[1]), .B1(N117), 
        .Y(N979) );
  AOI22X1TF U448 ( .A0(SUM_AB[8]), .A1(N82), .B0(N998), .B1(N1015), .Y(N999)
         );
  AOI22X1TF U449 ( .A0(DIVISION_HEAD[8]), .A1(N139), .B0(ZTEMP[8]), .B1(N116), 
        .Y(N1000) );
  INVX2TF U450 ( .A(N882), .Y(N210) );
  AOI31X1TF U451 ( .A0(N836), .A1(N835), .A2(N834), .B0(N924), .Y(N838) );
  AOI32X1TF U452 ( .A0(N833), .A1(OPER_B[2]), .A2(N922), .B0(N921), .B1(
        OPER_B[2]), .Y(N834) );
  AOI22X1TF U453 ( .A0(N920), .A1(OPER_B[3]), .B0(OPER_A[2]), .B1(N832), .Y(
        N835) );
  AOI31X1TF U454 ( .A0(N922), .A1(N156), .A2(N828), .B0(N827), .Y(N836) );
  OAI211X1TF U455 ( .A0(N1010), .A1(N1003), .B0(N1002), .C0(N1001), .Y(N660)
         );
  AOI22X1TF U456 ( .A0(DIVISION_HEAD[9]), .A1(N1012), .B0(ZTEMP[9]), .B1(N117), 
        .Y(N1002) );
  AOI211X1TF U457 ( .A0(N218), .A1(OPER_B[10]), .B0(N927), .C0(N928), .Y(N216)
         );
  AOI21X1TF U458 ( .A0(N975), .A1(N971), .B0(N910), .Y(N928) );
  AOI21X1TF U459 ( .A0(N926), .A1(N925), .B0(N924), .Y(N927) );
  AOI32X1TF U460 ( .A0(N923), .A1(OPER_B[10]), .A2(N922), .B0(N921), .B1(
        OPER_B[10]), .Y(N925) );
  AOI211X1TF U461 ( .A0(N920), .A1(OPER_B[11]), .B0(N919), .C0(N918), .Y(N926)
         );
  AOI21X1TF U462 ( .A0(N913), .A1(N917), .B0(N912), .Y(N914) );
  NOR3X1TF U463 ( .A(N911), .B(OPER_B[10]), .C(N923), .Y(N919) );
  AOI211X1TF U464 ( .A0(OPER_B[6]), .A1(N879), .B0(N878), .C0(N877), .Y(N880)
         );
  AOI21X1TF U465 ( .A0(N913), .A1(N876), .B0(N912), .Y(N874) );
  OAI31X1TF U466 ( .A0(N911), .A1(OPER_B[6]), .A2(N873), .B0(N872), .Y(N878)
         );
  AOI21X1TF U467 ( .A0(OPER_B[7]), .A1(N871), .B0(N870), .Y(N872) );
  OAI21X1TF U468 ( .A0(N911), .A1(N869), .B0(N868), .Y(N879) );
  AOI32X1TF U469 ( .A0(N394), .A1(N393), .A2(N392), .B0(N476), .B1(N393), .Y(
        N719) );
  OAI211X1TF U470 ( .A0(N390), .A1(N559), .B0(N389), .C0(N388), .Y(N391) );
  AOI22X1TF U471 ( .A0(X_IN[6]), .A1(N132), .B0(X_IN[5]), .B1(N100), .Y(N388)
         );
  AOI22X1TF U472 ( .A0(DIVISION_HEAD[3]), .A1(N735), .B0(SUM_AB[0]), .B1(N382), 
        .Y(N394) );
  OAI22X1TF U473 ( .A0(N476), .A1(N475), .B0(N474), .B1(N176), .Y(N711) );
  AOI211X1TF U474 ( .A0(N998), .A1(N494), .B0(N471), .C0(N470), .Y(N475) );
  OAI211X1TF U475 ( .A0(N469), .A1(N609), .B0(N468), .C0(N467), .Y(N470) );
  AOI22X1TF U476 ( .A0(XTEMP[9]), .A1(N89), .B0(N799), .B1(SUM_AB[12]), .Y(
        N467) );
  NOR2X1TF U477 ( .A(DIVISION_HEAD[12]), .B(N473), .Y(N466) );
  AOI22X1TF U478 ( .A0(X_IN[8]), .A1(N465), .B0(INTADD_0_N1), .B1(N489), .Y(
        N473) );
  OAI22X1TF U479 ( .A0(N143), .A1(N94), .B0(N464), .B1(N96), .Y(N471) );
  AOI32X1TF U480 ( .A0(N403), .A1(N461), .A2(N402), .B0(N476), .B1(N141), .Y(
        N718) );
  AOI211X1TF U481 ( .A0(N494), .A1(N977), .B0(N401), .C0(N400), .Y(N402) );
  OAI211X1TF U482 ( .A0(N559), .A1(N433), .B0(N399), .C0(N398), .Y(N400) );
  AOI21X1TF U483 ( .A0(DIVISION_HEAD[4]), .A1(N735), .B0(N397), .Y(N398) );
  OAI22X1TF U484 ( .A0(N141), .A1(N455), .B0(N749), .B1(N609), .Y(N397) );
  AOI22X1TF U485 ( .A0(DIVISION_HEAD[6]), .A1(N89), .B0(X_IN[7]), .B1(N131), 
        .Y(N399) );
  OAI22X1TF U486 ( .A0(N464), .A1(N396), .B0(N489), .B1(N748), .Y(N401) );
  AOI32X1TF U487 ( .A0(N432), .A1(N461), .A2(N431), .B0(N476), .B1(N151), .Y(
        N715) );
  AOI211X1TF U488 ( .A0(N494), .A1(N986), .B0(N430), .C0(N429), .Y(N431) );
  AOI22X1TF U489 ( .A0(DIVISION_HEAD[9]), .A1(N89), .B0(X_IN[9]), .B1(N100), 
        .Y(N427) );
  OAI22X1TF U490 ( .A0(N144), .A1(N94), .B0(N151), .B1(N455), .Y(N430) );
  OAI21X1TF U491 ( .A0(N451), .A1(N450), .B0(N461), .Y(N452) );
  AOI22X1TF U492 ( .A0(DIVISION_HEAD[11]), .A1(N89), .B0(X_IN[12]), .B1(N132), 
        .Y(N446) );
  AOI22X1TF U493 ( .A0(SUM_AB[6]), .A1(N127), .B0(N494), .B1(N992), .Y(N448)
         );
  OAI22X1TF U494 ( .A0(N145), .A1(N94), .B0(N443), .B1(N96), .Y(N451) );
  AOI22X1TF U495 ( .A0(SUM_AB[10]), .A1(N83), .B0(N1004), .B1(N1015), .Y(N1005) );
  AOI22X1TF U496 ( .A0(DIVISION_HEAD[10]), .A1(N139), .B0(ZTEMP[10]), .B1(N117), .Y(N1006) );
  OAI22X1TF U497 ( .A0(N514), .A1(N497), .B0(N496), .B1(N147), .Y(N709) );
  AOI21X1TF U498 ( .A0(N494), .A1(N1004), .B0(N493), .Y(N497) );
  OAI211X1TF U499 ( .A0(N501), .A1(N609), .B0(N492), .C0(N491), .Y(N493) );
  AOI22X1TF U500 ( .A0(XTEMP[11]), .A1(N89), .B0(SUM_AB[10]), .B1(N127), .Y(
        N492) );
  AOI32X1TF U501 ( .A0(N413), .A1(N461), .A2(N412), .B0(N476), .B1(N152), .Y(
        N717) );
  AOI211X1TF U502 ( .A0(DIVISION_HEAD[7]), .A1(N89), .B0(N411), .C0(N410), .Y(
        N412) );
  OAI211X1TF U503 ( .A0(N96), .A1(N749), .B0(N409), .C0(N408), .Y(N410) );
  AOI21X1TF U504 ( .A0(N494), .A1(N980), .B0(N407), .Y(N408) );
  OAI22X1TF U505 ( .A0(N141), .A1(N93), .B0(N152), .B1(N455), .Y(N407) );
  AOI22X1TF U506 ( .A0(X_IN[1]), .A1(N445), .B0(N799), .B1(SUM_AB[6]), .Y(N409) );
  OAI21X1TF U507 ( .A0(N501), .A1(N748), .B0(N404), .Y(N411) );
  AOI22X1TF U508 ( .A0(X_IN[8]), .A1(N132), .B0(X_IN[7]), .B1(N100), .Y(N404)
         );
  OAI211X1TF U509 ( .A0(N1010), .A1(N1009), .B0(N1008), .C0(N1007), .Y(N658)
         );
  AOI22X1TF U510 ( .A0(DIVISION_HEAD[11]), .A1(N139), .B0(ZTEMP[11]), .B1(N117), .Y(N1008) );
  OAI21X1TF U511 ( .A0(N760), .A1(N179), .B0(N563), .Y(N705) );
  OAI22X1TF U512 ( .A0(N562), .A1(N561), .B0(N762), .B1(N779), .Y(N563) );
  AOI22X1TF U513 ( .A0(Y_IN[0]), .A1(N790), .B0(DIVISION_REMA[1]), .B1(N113), 
        .Y(N560) );
  AOI21X1TF U514 ( .A0(N112), .A1(N650), .B0(N976), .Y(N562) );
  INVX2TF U515 ( .A(SUM_AB[0]), .Y(N976) );
  INVX2TF U516 ( .A(N922), .Y(N911) );
  OAI211X1TF U517 ( .A0(N1019), .A1(N1018), .B0(N1017), .C0(N1016), .Y(N657)
         );
  AOI32X1TF U518 ( .A0(N1018), .A1(N1015), .A2(N1014), .B0(N1013), .B1(N1015), 
        .Y(N1016) );
  AOI211X4TF U519 ( .A0(N975), .A1(N974), .B0(N973), .C0(N116), .Y(N1015) );
  INVX2TF U520 ( .A(N969), .Y(N973) );
  AOI22X1TF U521 ( .A0(DIVISION_HEAD[12]), .A1(N139), .B0(ZTEMP[12]), .B1(N117), .Y(N1017) );
  OAI31X1TF U522 ( .A0(N967), .A1(N56), .A2(N971), .B0(N966), .Y(N968) );
  AOI31X1TF U523 ( .A0(N178), .A1(N56), .A2(N965), .B0(N964), .Y(N966) );
  AOI31X1TF U524 ( .A0(N960), .A1(N959), .A2(N958), .B0(N957), .Y(N963) );
  OAI31X1TF U525 ( .A0(N956), .A1(N955), .A2(N954), .B0(N953), .Y(N957) );
  OAI22X1TF U526 ( .A0(N514), .A1(N359), .B0(N358), .B1(N171), .Y(N723) );
  AOI211X1TF U527 ( .A0(N494), .A1(N1013), .B0(N356), .C0(N355), .Y(N359) );
  OAI31X1TF U528 ( .A0(XTEMP[12]), .A1(N357), .A2(N510), .B0(N354), .Y(N355)
         );
  OAI22X1TF U529 ( .A0(N112), .A1(N1018), .B0(N503), .B1(N96), .Y(N356) );
  OAI22X1TF U530 ( .A0(N192), .A1(N752), .B0(N760), .B1(N174), .Y(N688) );
  AOI211X1TF U531 ( .A0(N992), .A1(N796), .B0(N751), .C0(N750), .Y(N752) );
  OAI211X1TF U532 ( .A0(N749), .A1(N748), .B0(N756), .C0(N747), .Y(N750) );
  AOI22X1TF U533 ( .A0(DIVISION_REMA[7]), .A1(N113), .B0(SUM_AB[6]), .B1(N137), 
        .Y(N747) );
  OAI21X1TF U534 ( .A0(N201), .A1(N96), .B0(N745), .Y(N751) );
  AOI22X1TF U535 ( .A0(Y_IN[6]), .A1(N790), .B0(DIVISION_REMA[5]), .B1(N735), 
        .Y(N745) );
  AOI21X1TF U536 ( .A0(SUM_AB[6]), .A1(N444), .B0(N454), .Y(N992) );
  OAI22X1TF U537 ( .A0(N514), .A1(N513), .B0(N512), .B1(N155), .Y(N708) );
  OAI21X1TF U538 ( .A0(N508), .A1(N1009), .B0(N507), .Y(N509) );
  AOI211X1TF U539 ( .A0(SUM_AB[11]), .A1(N127), .B0(N505), .C0(N504), .Y(N507)
         );
  OAI22X1TF U540 ( .A0(N147), .A1(N93), .B0(N501), .B1(N95), .Y(N505) );
  OAI22X1TF U541 ( .A0(N514), .A1(N486), .B0(N485), .B1(N529), .Y(N710) );
  AOI211X1TF U542 ( .A0(SUM_AB[9]), .A1(N130), .B0(N483), .C0(N482), .Y(N486)
         );
  OAI211X1TF U543 ( .A0(N1003), .A1(N508), .B0(N481), .C0(N480), .Y(N482) );
  INVX2TF U544 ( .A(INTADD_0_N1), .Y(N465) );
  OAI22X1TF U545 ( .A0(N176), .A1(N94), .B0(N489), .B1(N609), .Y(N483) );
  AOI32X1TF U546 ( .A0(N798), .A1(N815), .A2(N797), .B0(N813), .B1(N173), .Y(
        N684) );
  AOI21X1TF U547 ( .A0(N796), .A1(N1004), .B0(N795), .Y(N797) );
  AOI22X1TF U548 ( .A0(X_IN[2]), .A1(N100), .B0(X_IN[4]), .B1(N806), .Y(N791)
         );
  AOI22X1TF U549 ( .A0(DIVISION_HEAD[0]), .A1(N126), .B0(DIVISION_HEAD[1]), 
        .B1(N805), .Y(N792) );
  AOI22X1TF U550 ( .A0(Y_IN[10]), .A1(N790), .B0(X_IN[3]), .B1(N132), .Y(N793)
         );
  AOI21X1TF U551 ( .A0(SUM_AB[10]), .A1(N487), .B0(N500), .Y(N1004) );
  AOI22X1TF U552 ( .A0(N799), .A1(SUM_AB[1]), .B0(SUM_AB[10]), .B1(N138), .Y(
        N798) );
  AOI32X1TF U553 ( .A0(N462), .A1(N461), .A2(N460), .B0(N476), .B1(N143), .Y(
        N712) );
  OAI211X1TF U554 ( .A0(N508), .A1(N997), .B0(N457), .C0(N456), .Y(N458) );
  AOI22X1TF U555 ( .A0(DIVISION_HEAD[12]), .A1(N88), .B0(X_IN[12]), .B1(N99), 
        .Y(N456) );
  AOI22X1TF U556 ( .A0(DIVISION_HEAD[11]), .A1(N805), .B0(DIVISION_HEAD[10]), 
        .B1(N126), .Y(N457) );
  OAI22X1TF U557 ( .A0(N464), .A1(N609), .B0(N559), .B1(N499), .Y(N459) );
  OAI21X1TF U558 ( .A0(N813), .A1(N556), .B0(N555), .Y(N706) );
  OAI21X1TF U559 ( .A0(N813), .A1(N805), .B0(DIVISION_HEAD[3]), .Y(N555) );
  AOI211X1TF U560 ( .A0(DIVISION_HEAD[2]), .A1(N126), .B0(N554), .C0(N553), 
        .Y(N556) );
  AOI22X1TF U561 ( .A0(N799), .A1(SUM_AB[3]), .B0(N1013), .B1(N796), .Y(N550)
         );
  NOR2X1TF U562 ( .A(N1018), .B(N1014), .Y(N1013) );
  AOI22X1TF U563 ( .A0(N941), .A1(SUM_AB[12]), .B0(X_IN[5]), .B1(N132), .Y(
        N551) );
  AOI22X1TF U564 ( .A0(X_IN[4]), .A1(N100), .B0(X_IN[6]), .B1(N806), .Y(N552)
         );
  OAI22X1TF U565 ( .A0(N549), .A1(N803), .B0(N548), .B1(N96), .Y(N554) );
  OAI22X1TF U566 ( .A0(N192), .A1(N654), .B0(N760), .B1(N159), .Y(N693) );
  AOI21X1TF U567 ( .A0(SUM_AB[1]), .A1(N138), .B0(N653), .Y(N654) );
  AOI22X1TF U568 ( .A0(DIVISION_REMA[0]), .A1(N735), .B0(N796), .B1(N977), .Y(
        N651) );
  AOI21X1TF U569 ( .A0(SUM_AB[1]), .A1(SUM_AB[0]), .B0(N405), .Y(N977) );
  AOI22X1TF U570 ( .A0(Y_IN[1]), .A1(N790), .B0(DIVISION_REMA[2]), .B1(N114), 
        .Y(N652) );
  AOI22X1TF U571 ( .A0(N192), .A1(N146), .B0(N780), .B1(N779), .Y(N686) );
  AOI211X1TF U572 ( .A0(DIVISION_REMA[7]), .A1(N735), .B0(N778), .C0(N777), 
        .Y(N780) );
  OAI211X1TF U573 ( .A0(N169), .A1(N776), .B0(N775), .C0(N774), .Y(N777) );
  AOI22X1TF U574 ( .A0(N773), .A1(N772), .B0(N998), .B1(N796), .Y(N774) );
  AOI21X1TF U575 ( .A0(SUM_AB[8]), .A1(N463), .B0(N478), .Y(N998) );
  AOI32X1TF U576 ( .A0(N771), .A1(N770), .A2(N769), .B0(N768), .B1(N770), .Y(
        N772) );
  OAI32X1TF U577 ( .A0(N767), .A1(N766), .A2(X_IN[0]), .B0(N765), .B1(N767), 
        .Y(N770) );
  AOI22X1TF U578 ( .A0(DIVISION_REMA[8]), .A1(N762), .B0(SUM_AB[8]), .B1(N137), 
        .Y(N775) );
  OAI21X1TF U579 ( .A0(N176), .A1(N98), .B0(N239), .Y(FOUT[8]) );
  AOI21X1TF U580 ( .A0(N220), .A1(DIVISION_REMA[8]), .B0(N238), .Y(N239) );
  OAI22X1TF U581 ( .A0(N173), .A1(N81), .B0(N147), .B1(N86), .Y(N238) );
  AOI22X1TF U582 ( .A0(N476), .A1(N145), .B0(N442), .B1(N461), .Y(N714) );
  AOI21X1TF U583 ( .A0(DIVISION_HEAD[8]), .A1(N126), .B0(N435), .Y(N436) );
  OAI22X1TF U584 ( .A0(N145), .A1(N455), .B0(N508), .B1(N991), .Y(N435) );
  AOI22X1TF U585 ( .A0(DIVISION_HEAD[10]), .A1(N88), .B0(X_IN[10]), .B1(N99), 
        .Y(N438) );
  OAI22X1TF U586 ( .A0(N443), .A1(N609), .B0(N559), .B1(N477), .Y(N441) );
  OAI22X1TF U587 ( .A0(N192), .A1(N740), .B0(N760), .B1(N170), .Y(N690) );
  AOI211X1TF U588 ( .A0(SUM_AB[4]), .A1(N138), .B0(N739), .C0(N738), .Y(N740)
         );
  OAI211X1TF U589 ( .A0(N737), .A1(N96), .B0(N756), .C0(N736), .Y(N738) );
  AOI22X1TF U590 ( .A0(DIVISION_REMA[5]), .A1(N114), .B0(N796), .B1(N986), .Y(
        N736) );
  AOI21X1TF U591 ( .A0(SUM_AB[4]), .A1(N424), .B0(N434), .Y(N986) );
  OAI22X1TF U592 ( .A0(N201), .A1(N803), .B0(N166), .B1(N94), .Y(N739) );
  OAI22X1TF U593 ( .A0(N192), .A1(N729), .B0(N760), .B1(N172), .Y(N692) );
  AOI211X1TF U594 ( .A0(SUM_AB[2]), .A1(N138), .B0(N728), .C0(N727), .Y(N729)
         );
  OAI211X1TF U595 ( .A0(N656), .A1(N96), .B0(N756), .C0(N655), .Y(N727) );
  AOI22X1TF U596 ( .A0(DIVISION_REMA[3]), .A1(N114), .B0(N796), .B1(N980), .Y(
        N655) );
  AOI21X1TF U597 ( .A0(SUM_AB[2]), .A1(N406), .B0(N416), .Y(N980) );
  NOR2X1TF U598 ( .A(SUM_AB[0]), .B(SUM_AB[1]), .Y(N405) );
  OAI22X1TF U599 ( .A0(N737), .A1(N803), .B0(N159), .B1(N94), .Y(N728) );
  OAI21X1TF U600 ( .A0(N151), .A1(N98), .B0(N231), .Y(FOUT[4]) );
  AOI21X1TF U601 ( .A0(N220), .A1(DIVISION_REMA[4]), .B0(N230), .Y(N231) );
  OAI22X1TF U602 ( .A0(N154), .A1(N87), .B0(N174), .B1(N81), .Y(N230) );
  AOI32X1TF U603 ( .A0(N423), .A1(N461), .A2(N422), .B0(N476), .B1(N144), .Y(
        N716) );
  AOI211X1TF U604 ( .A0(DIVISION_HEAD[8]), .A1(N89), .B0(N421), .C0(N420), .Y(
        N422) );
  OAI211X1TF U605 ( .A0(N559), .A1(N453), .B0(N419), .C0(N418), .Y(N420) );
  AOI21X1TF U606 ( .A0(DIVISION_HEAD[6]), .A1(N735), .B0(N417), .Y(N418) );
  OAI22X1TF U607 ( .A0(N144), .A1(N455), .B0(N508), .B1(N985), .Y(N417) );
  INVX2TF U608 ( .A(N494), .Y(N508) );
  NOR2X2TF U609 ( .A(N395), .B(N1018), .Y(N494) );
  AOI22X1TF U610 ( .A0(X_IN[2]), .A1(N445), .B0(X_IN[1]), .B1(N801), .Y(N419)
         );
  INVX2TF U611 ( .A(N609), .Y(N445) );
  NAND2X2TF U612 ( .A(MODE_TYPE[1]), .B(N353), .Y(N609) );
  OAI21X1TF U613 ( .A0(N503), .A1(N748), .B0(N414), .Y(N421) );
  AOI22X1TF U614 ( .A0(X_IN[8]), .A1(N100), .B0(X_IN[9]), .B1(N132), .Y(N414)
         );
  INVX2TF U615 ( .A(N806), .Y(N748) );
  AOI31X1TF U616 ( .A0(N941), .A1(N73), .A2(N564), .B0(N350), .Y(N386) );
  OAI211X1TF U617 ( .A0(N73), .A1(N376), .B0(N360), .C0(N349), .Y(N350) );
  OAI211X1TF U618 ( .A0(N960), .A1(N348), .B0(N567), .C0(N601), .Y(N349) );
  NOR2X1TF U619 ( .A(N372), .B(N944), .Y(N360) );
  INVX2TF U620 ( .A(N395), .Y(N372) );
  INVX2TF U621 ( .A(N618), .Y(N376) );
  NOR2X1TF U622 ( .A(N153), .B(N749), .Y(INTADD_0_CI) );
  INVX2TF U623 ( .A(X_IN[0]), .Y(N749) );
  NOR2X1TF U624 ( .A(PRE_WORK), .B(N365), .Y(N603) );
  INVX2TF U625 ( .A(N600), .Y(N567) );
  OAI211X1TF U626 ( .A0(N856), .A1(N855), .B0(N854), .C0(N853), .Y(N678) );
  AOI32X1TF U627 ( .A0(N937), .A1(OPER_B[4]), .A2(N852), .B0(N884), .B1(
        OPER_B[4]), .Y(N853) );
  AOI211X1TF U628 ( .A0(N858), .A1(OPER_B[5]), .B0(N851), .C0(N850), .Y(N854)
         );
  OAI31X1TF U629 ( .A0(N934), .A1(OPER_A[4]), .A2(N849), .B0(N205), .Y(N850)
         );
  AOI21X1TF U630 ( .A0(N106), .A1(C152_DATA4_4), .B0(N207), .Y(N205) );
  NOR3X1TF U631 ( .A(OPER_B[4]), .B(N852), .C(N109), .Y(N851) );
  AOI21X1TF U632 ( .A0(N931), .A1(N849), .B0(N848), .Y(N855) );
  INVX2TF U633 ( .A(N932), .Y(N848) );
  AOI211X1TF U634 ( .A0(N107), .A1(C152_DATA4_5), .B0(N860), .C0(N211), .Y(
        N212) );
  OAI31X1TF U635 ( .A0(OPER_B[5]), .A1(N859), .A2(N109), .B0(N905), .Y(N860)
         );
  OAI211X1TF U636 ( .A0(SIGN_Y), .A1(N965), .B0(N221), .C0(N971), .Y(N905) );
  AOI22X1TF U637 ( .A0(N858), .A1(OPER_B[6]), .B0(N857), .B1(N862), .Y(N867)
         );
  NOR2X1TF U638 ( .A(N934), .B(OPER_A[5]), .Y(N857) );
  INVX2TF U639 ( .A(N894), .Y(N858) );
  AOI22X1TF U640 ( .A0(OPER_B[5]), .A1(N864), .B0(OPER_A[5]), .B1(N863), .Y(
        N866) );
  OAI21X1TF U641 ( .A0(N934), .A1(N862), .B0(N932), .Y(N863) );
  OAI21X1TF U642 ( .A0(N109), .A1(N861), .B0(N935), .Y(N864) );
  OAI21X1TF U643 ( .A0(N141), .A1(N97), .B0(N225), .Y(FOUT[1]) );
  AOI21X1TF U644 ( .A0(N220), .A1(DIVISION_REMA[1]), .B0(N224), .Y(N225) );
  OAI22X1TF U645 ( .A0(N144), .A1(N86), .B0(N166), .B1(N80), .Y(N224) );
  OAI211X1TF U646 ( .A0(N894), .A1(N160), .B0(N893), .C0(N892), .Y(N675) );
  AOI211X1TF U647 ( .A0(OPER_A[7]), .A1(N890), .B0(N889), .C0(N888), .Y(N893)
         );
  INVX2TF U648 ( .A(N208), .Y(N888) );
  AOI211X1TF U649 ( .A0(N106), .A1(C152_DATA4_7), .B0(N207), .C0(N206), .Y(
        N208) );
  NOR3X1TF U650 ( .A(N108), .B(OPER_B[7]), .C(N887), .Y(N206) );
  OR2X2TF U651 ( .A(N930), .B(N886), .Y(N207) );
  NOR2X1TF U652 ( .A(N967), .B(N830), .Y(N870) );
  INVX2TF U653 ( .A(N885), .Y(N889) );
  AOI32X1TF U654 ( .A0(OPER_B[7]), .A1(N937), .A2(N887), .B0(N884), .B1(
        OPER_B[7]), .Y(N885) );
  INVX2TF U655 ( .A(N935), .Y(N884) );
  OAI21X1TF U656 ( .A0(N934), .A1(N891), .B0(N932), .Y(N890) );
  NOR3X1TF U657 ( .A(N73), .B(N178), .C(N965), .Y(N964) );
  OAI22X1TF U658 ( .A0(N190), .A1(N201), .B0(N202), .B1(OFFSET[2]), .Y(C2_Z_4)
         );
  INVX2TF U659 ( .A(Y_IN[4]), .Y(N201) );
  OAI22X1TF U660 ( .A0(N190), .A1(N200), .B0(N202), .B1(OFFSET[3]), .Y(C2_Z_5)
         );
  OAI22X1TF U661 ( .A0(N190), .A1(N199), .B0(N202), .B1(OFFSET[4]), .Y(C2_Z_6)
         );
  OAI22X1TF U662 ( .A0(N190), .A1(N194), .B0(N202), .B1(OFFSET[5]), .Y(C2_Z_7)
         );
  OAI22X1TF U663 ( .A0(N190), .A1(N761), .B0(N202), .B1(OFFSET[6]), .Y(C2_Z_8)
         );
  OAI22X1TF U664 ( .A0(N190), .A1(N783), .B0(N202), .B1(OFFSET[7]), .Y(C2_Z_9)
         );
  OAI22X1TF U665 ( .A0(N190), .A1(N548), .B0(N133), .B1(OFFSET[8]), .Y(C2_Z_10) );
  OAI22X1TF U666 ( .A0(N190), .A1(N804), .B0(N133), .B1(OFFSET[9]), .Y(C2_Z_11) );
  NOR2X1TF U667 ( .A(OPER_B[9]), .B(N908), .Y(N923) );
  NOR2X1TF U668 ( .A(N869), .B(OPER_B[6]), .Y(N887) );
  INVX2TF U669 ( .A(N873), .Y(N869) );
  NOR2X1TF U670 ( .A(OPER_B[5]), .B(N861), .Y(N873) );
  NOR2X1TF U671 ( .A(OPER_B[3]), .B(N841), .Y(N852) );
  AOI211X1TF U672 ( .A0(N56), .A1(N965), .B0(SIGN_Y), .C0(N910), .Y(N930) );
  NOR2X1TF U673 ( .A(OPER_A[9]), .B(N909), .Y(N917) );
  NOR2X1TF U674 ( .A(OPER_A[7]), .B(N891), .Y(N898) );
  NOR2X1TF U675 ( .A(OPER_A[5]), .B(N862), .Y(N876) );
  NOR2X1TF U676 ( .A(OPER_A[3]), .B(N840), .Y(N849) );
  OAI211X1TF U677 ( .A0(N177), .A1(N938), .B0(N847), .C0(N846), .Y(N679) );
  AOI211X1TF U678 ( .A0(OPER_A[3]), .A1(N845), .B0(N844), .C0(N843), .Y(N846)
         );
  OAI31X1TF U679 ( .A0(N934), .A1(OPER_A[3]), .A2(N842), .B0(N204), .Y(N843)
         );
  AOI21X1TF U680 ( .A0(C152_DATA4_3), .A1(N106), .B0(N906), .Y(N204) );
  OAI22X1TF U681 ( .A0(N970), .A1(N730), .B0(N202), .B1(OFFSET[1]), .Y(C2_Z_3)
         );
  INVX2TF U682 ( .A(DP_OP_333_124_4748_N57), .Y(N202) );
  OAI32X1TF U683 ( .A0(N183), .A1(N108), .A2(N841), .B0(N935), .B1(N183), .Y(
        N844) );
  INVX2TF U684 ( .A(N868), .Y(N921) );
  AOI32X1TF U685 ( .A0(N606), .A1(N347), .A2(N823), .B0(N946), .B1(N346), .Y(
        N868) );
  INVX2TF U686 ( .A(N940), .Y(N946) );
  OAI21X1TF U687 ( .A0(N934), .A1(N840), .B0(N932), .Y(N845) );
  INVX2TF U688 ( .A(N831), .Y(N912) );
  AOI21X1TF U689 ( .A0(N565), .A1(N346), .B0(N564), .Y(N831) );
  INVX2TF U690 ( .A(N842), .Y(N840) );
  NOR3X1TF U691 ( .A(OPER_A[2]), .B(OPER_A[1]), .C(OPER_A[0]), .Y(N842) );
  INVX2TF U692 ( .A(N931), .Y(N934) );
  NOR2X2TF U693 ( .A(N924), .B(N916), .Y(N931) );
  INVX2TF U694 ( .A(N904), .Y(N924) );
  AOI31X1TF U695 ( .A0(N937), .A1(N183), .A2(N841), .B0(N882), .Y(N847) );
  OAI21X1TF U696 ( .A0(N975), .A1(N910), .B0(N837), .Y(N882) );
  INVX2TF U697 ( .A(N910), .Y(N221) );
  INVX2TF U698 ( .A(N345), .Y(N959) );
  INVX2TF U699 ( .A(N566), .Y(N949) );
  NOR2X1TF U700 ( .A(OPER_B[1]), .B(OPER_B[0]), .Y(N833) );
  INVX2TF U701 ( .A(N346), .Y(N347) );
  INVX2TF U702 ( .A(N606), .Y(N822) );
  NOR2X2TF U703 ( .A(N604), .B(N632), .Y(N823) );
  AOI221X1TF U704 ( .A0(N128), .A1(N158), .B0(N181), .B1(N91), .C0(N818), .Y(
        N819) );
  AOI22X1TF U705 ( .A0(\INDEX[2] ), .A1(N90), .B0(N124), .B1(\RSHT_BITS[3] ), 
        .Y(N817) );
  AOI32X1TF U706 ( .A0(N940), .A1(N953), .A2(N369), .B0(N955), .B1(N953), .Y(
        N343) );
  OR2X2TF U707 ( .A(N632), .B(N149), .Y(N369) );
  INVX2TF U708 ( .A(N604), .Y(N643) );
  OAI21X1TF U709 ( .A0(N345), .A1(N939), .B0(N341), .Y(N608) );
  OAI21X1TF U710 ( .A0(N571), .A1(N565), .B0(N342), .Y(N341) );
  NOR2X2TF U711 ( .A(\RSHT_BITS[3] ), .B(N592), .Y(N606) );
  NOR3X1TF U712 ( .A(N121), .B(N122), .C(N954), .Y(N821) );
  INVX2TF U713 ( .A(N960), .Y(N967) );
  NOR2X1TF U714 ( .A(SIGN_Y), .B(N110), .Y(N907) );
  OAI22X1TF U715 ( .A0(Y_IN[12]), .A1(N176), .B0(N337), .B1(N336), .Y(N338) );
  OAI31X1TF U716 ( .A0(N335), .A1(DIVISION_HEAD[10]), .A2(N548), .B0(N334), 
        .Y(N336) );
  AOI22X1TF U717 ( .A0(Y_IN[11]), .A1(N143), .B0(N333), .B1(N332), .Y(N334) );
  OAI22X1TF U718 ( .A0(DIVISION_HEAD[8]), .A1(N761), .B0(DIVISION_HEAD[9]), 
        .B1(N783), .Y(N332) );
  INVX2TF U719 ( .A(N331), .Y(N333) );
  NOR2X1TF U720 ( .A(Y_IN[11]), .B(N143), .Y(N335) );
  AOI211X1TF U721 ( .A0(DIVISION_HEAD[8]), .A1(N761), .B0(N330), .C0(N331), 
        .Y(N337) );
  OAI21X1TF U722 ( .A0(Y_IN[11]), .A1(N143), .B0(N329), .Y(N331) );
  AOI22X1TF U723 ( .A0(DIVISION_HEAD[10]), .A1(N548), .B0(DIVISION_HEAD[9]), 
        .B1(N783), .Y(N329) );
  AOI21X1TF U724 ( .A0(N84), .A1(N144), .B0(N328), .Y(N330) );
  AOI211X1TF U725 ( .A0(N327), .A1(DIVISION_HEAD[6]), .B0(N326), .C0(N325), 
        .Y(N328) );
  NOR2X1TF U726 ( .A(N84), .B(N144), .Y(N326) );
  AOI21X1TF U727 ( .A0(N193), .A1(N141), .B0(N324), .Y(N327) );
  AOI211X1TF U728 ( .A0(N323), .A1(DIVISION_HEAD[4]), .B0(N322), .C0(N321), 
        .Y(N324) );
  NOR2X1TF U729 ( .A(Y_IN[5]), .B(N141), .Y(N322) );
  AOI21X1TF U730 ( .A0(Y_IN[3]), .A1(N148), .B0(N320), .Y(N323) );
  OAI32X1TF U731 ( .A0(N319), .A1(DIVISION_HEAD[2]), .A2(N737), .B0(N318), 
        .B1(N319), .Y(N320) );
  OAI211X1TF U732 ( .A0(Y_IN[2]), .A1(N163), .B0(N317), .C0(N316), .Y(N318) );
  NOR2X1TF U733 ( .A(Y_IN[3]), .B(N148), .Y(N319) );
  INVX2TF U734 ( .A(Y_IN[12]), .Y(N549) );
  OAI21X1TF U735 ( .A0(N144), .A1(N97), .B0(N229), .Y(FOUT[3]) );
  AOI21X1TF U736 ( .A0(N220), .A1(DIVISION_REMA[3]), .B0(N228), .Y(N229) );
  OAI22X1TF U737 ( .A0(N145), .A1(N86), .B0(N167), .B1(N80), .Y(N228) );
  OAI21X1TF U738 ( .A0(N143), .A1(N98), .B0(N237), .Y(FOUT[7]) );
  AOI21X1TF U739 ( .A0(N220), .A1(DIVISION_REMA[7]), .B0(N236), .Y(N237) );
  OAI22X1TF U740 ( .A0(N169), .A1(N81), .B0(N529), .B1(N87), .Y(N236) );
  OAI21X1TF U741 ( .A0(N145), .A1(N97), .B0(N233), .Y(FOUT[5]) );
  AOI21X1TF U742 ( .A0(N220), .A1(DIVISION_REMA[5]), .B0(N232), .Y(N233) );
  OAI22X1TF U743 ( .A0(N143), .A1(N86), .B0(N168), .B1(N80), .Y(N232) );
  OAI21X1TF U744 ( .A0(N152), .A1(N97), .B0(N227), .Y(FOUT[2]) );
  AOI21X1TF U745 ( .A0(N220), .A1(DIVISION_REMA[2]), .B0(N226), .Y(N227) );
  OAI22X1TF U746 ( .A0(N151), .A1(N86), .B0(N170), .B1(N80), .Y(N226) );
  OAI21X1TF U747 ( .A0(N154), .A1(N98), .B0(N235), .Y(FOUT[6]) );
  AOI21X1TF U748 ( .A0(N220), .A1(DIVISION_REMA[6]), .B0(N234), .Y(N235) );
  OAI22X1TF U749 ( .A0(N176), .A1(N87), .B0(N146), .B1(N80), .Y(N234) );
  OAI21X1TF U750 ( .A0(N760), .A1(N168), .B0(N759), .Y(N687) );
  OAI21X1TF U751 ( .A0(N758), .A1(N757), .B0(N779), .Y(N759) );
  INVX2TF U752 ( .A(N192), .Y(N779) );
  OAI211X1TF U753 ( .A0(N146), .A1(N776), .B0(N756), .C0(N755), .Y(N757) );
  AOI22X1TF U754 ( .A0(DIVISION_REMA[6]), .A1(N735), .B0(SUM_AB[7]), .B1(N137), 
        .Y(N755) );
  OAI211X1TF U755 ( .A0(N809), .A1(N997), .B0(N754), .C0(N753), .Y(N758) );
  AOI22X1TF U756 ( .A0(X_IN[1]), .A1(N806), .B0(X_IN[0]), .B1(N132), .Y(N753)
         );
  OAI21X1TF U757 ( .A0(N454), .A1(N453), .B0(N463), .Y(N997) );
  OAI22X1TF U758 ( .A0(N192), .A1(N734), .B0(N760), .B1(N166), .Y(N691) );
  AOI211X1TF U759 ( .A0(SUM_AB[3]), .A1(N138), .B0(N733), .C0(N732), .Y(N734)
         );
  OAI211X1TF U760 ( .A0(N809), .A1(N985), .B0(N756), .C0(N731), .Y(N732) );
  OAI21X1TF U761 ( .A0(N416), .A1(N415), .B0(N424), .Y(N985) );
  OAI22X1TF U762 ( .A0(N730), .A1(N803), .B0(N172), .B1(N94), .Y(N733) );
  OAI22X1TF U763 ( .A0(N192), .A1(N744), .B0(N760), .B1(N167), .Y(N689) );
  AOI211X1TF U764 ( .A0(SUM_AB[5]), .A1(N138), .B0(N743), .C0(N742), .Y(N744)
         );
  OAI211X1TF U765 ( .A0(N809), .A1(N991), .B0(N756), .C0(N741), .Y(N742) );
  AOI222X4TF U766 ( .A0(N766), .A1(N99), .B0(N764), .B1(N131), .C0(N558), .C1(
        N806), .Y(N756) );
  OAI21X1TF U767 ( .A0(N434), .A1(N433), .B0(N444), .Y(N991) );
  INVX2TF U768 ( .A(N803), .Y(N790) );
  NOR3X1TF U769 ( .A(N773), .B(N126), .C(N557), .Y(N781) );
  AOI32X1TF U770 ( .A0(N789), .A1(N815), .A2(N788), .B0(N813), .B1(N169), .Y(
        N685) );
  OAI211X1TF U771 ( .A0(N809), .A1(N1003), .B0(N785), .C0(N784), .Y(N786) );
  AOI22X1TF U772 ( .A0(DIVISION_HEAD[1]), .A1(N114), .B0(X_IN[1]), .B1(N99), 
        .Y(N784) );
  OAI21X1TF U773 ( .A0(N478), .A1(N477), .B0(N487), .Y(N1003) );
  OAI21X1TF U774 ( .A0(N783), .A1(N803), .B0(N782), .Y(N787) );
  AOI22X1TF U775 ( .A0(DIVISION_REMA[8]), .A1(N126), .B0(N799), .B1(SUM_AB[0]), 
        .Y(N782) );
  AOI22X1TF U776 ( .A0(DIVISION_HEAD[0]), .A1(N805), .B0(SUM_AB[9]), .B1(N138), 
        .Y(N789) );
  AOI32X1TF U777 ( .A0(N816), .A1(N815), .A2(N814), .B0(N813), .B1(N163), .Y(
        N683) );
  AOI211X1TF U778 ( .A0(DIVISION_HEAD[3]), .A1(N114), .B0(N811), .C0(N810), 
        .Y(N814) );
  OAI211X1TF U779 ( .A0(N809), .A1(N1009), .B0(N808), .C0(N807), .Y(N810) );
  AOI22X1TF U780 ( .A0(X_IN[3]), .A1(N99), .B0(X_IN[5]), .B1(N806), .Y(N807)
         );
  AND2X2TF U781 ( .A(N763), .B(N768), .Y(N765) );
  INVX2TF U782 ( .A(N387), .Y(N773) );
  AOI22X1TF U783 ( .A0(DIVISION_HEAD[1]), .A1(N126), .B0(DIVISION_HEAD[2]), 
        .B1(N805), .Y(N808) );
  INVX2TF U784 ( .A(N455), .Y(N805) );
  OAI21X1TF U785 ( .A0(N500), .A1(N499), .B0(N1014), .Y(N1009) );
  INVX2TF U786 ( .A(SUM_AB[11]), .Y(N499) );
  INVX2TF U787 ( .A(SUM_AB[9]), .Y(N477) );
  INVX2TF U788 ( .A(SUM_AB[7]), .Y(N453) );
  NOR2X1TF U789 ( .A(SUM_AB[6]), .B(N444), .Y(N454) );
  INVX2TF U790 ( .A(SUM_AB[5]), .Y(N433) );
  NOR2X1TF U791 ( .A(SUM_AB[4]), .B(N424), .Y(N434) );
  INVX2TF U792 ( .A(SUM_AB[3]), .Y(N415) );
  NOR3X1TF U793 ( .A(SUM_AB[0]), .B(SUM_AB[2]), .C(SUM_AB[1]), .Y(N416) );
  INVX2TF U794 ( .A(N796), .Y(N809) );
  NOR2X2TF U795 ( .A(N1018), .B(N650), .Y(N796) );
  INVX2TF U796 ( .A(SUM_AB[12]), .Y(N1018) );
  OAI21X1TF U797 ( .A0(N804), .A1(N803), .B0(N802), .Y(N811) );
  INVX2TF U798 ( .A(N95), .Y(N801) );
  NAND2X2TF U799 ( .A(N353), .B(N312), .Y(N803) );
  INVX2TF U800 ( .A(N813), .Y(N815) );
  AOI32X1TF U801 ( .A0(N120), .A1(N56), .A2(N564), .B0(N618), .B1(N73), .Y(
        N545) );
  INVX2TF U802 ( .A(N353), .Y(N640) );
  AOI31X1TF U803 ( .A0(N122), .A1(N385), .A2(N384), .B0(N383), .Y(N547) );
  INVX2TF U804 ( .A(N305), .Y(N764) );
  OAI211X1TF U805 ( .A0(X_IN[12]), .A1(N548), .B0(N304), .C0(N303), .Y(N305)
         );
  OAI22X1TF U806 ( .A0(Y_IN[10]), .A1(N302), .B0(N301), .B1(N300), .Y(N303) );
  OAI22X1TF U807 ( .A0(X_IN[10]), .A1(N299), .B0(X_IN[11]), .B1(N783), .Y(N300) );
  OAI21X1TF U808 ( .A0(Y_IN[9]), .A1(N298), .B0(Y_IN[8]), .Y(N299) );
  AOI211X1TF U809 ( .A0(X_IN[10]), .A1(N761), .B0(N297), .C0(N296), .Y(N301)
         );
  AOI21X1TF U810 ( .A0(Y_IN[7]), .A1(N501), .B0(N295), .Y(N296) );
  AOI211X1TF U811 ( .A0(X_IN[8]), .A1(N294), .B0(N293), .C0(N292), .Y(N295) );
  NOR2X1TF U812 ( .A(N84), .B(N501), .Y(N293) );
  AOI21X1TF U813 ( .A0(N193), .A1(N469), .B0(N291), .Y(N294) );
  AOI211X1TF U814 ( .A0(X_IN[6]), .A1(N290), .B0(N289), .C0(N288), .Y(N291) );
  NOR2X1TF U815 ( .A(N193), .B(N469), .Y(N289) );
  AOI32X1TF U816 ( .A0(N287), .A1(N286), .A2(N316), .B0(N285), .B1(N286), .Y(
        N290) );
  OAI22X1TF U817 ( .A0(X_IN[4]), .A1(N737), .B0(N101), .B1(N730), .Y(N285) );
  OAI32X1TF U818 ( .A0(N284), .A1(N85), .A2(N314), .B0(X_IN[2]), .B1(N284), 
        .Y(N287) );
  INVX2TF U819 ( .A(X_IN[7]), .Y(N469) );
  INVX2TF U820 ( .A(X_IN[9]), .Y(N501) );
  NOR2X1TF U821 ( .A(Y_IN[9]), .B(N298), .Y(N297) );
  INVX2TF U822 ( .A(X_IN[11]), .Y(N298) );
  NOR2X1TF U823 ( .A(Y_IN[12]), .B(Y_IN[11]), .Y(N304) );
  INVX2TF U824 ( .A(N769), .Y(N558) );
  OR2X2TF U825 ( .A(MODE_TYPE[0]), .B(N312), .Y(N768) );
  INVX2TF U826 ( .A(MODE_TYPE[1]), .Y(N312) );
  OAI31X1TF U827 ( .A0(N280), .A1(N279), .A2(N278), .B0(N277), .Y(N281) );
  INVX2TF U828 ( .A(Y_IN[11]), .Y(N804) );
  NOR2X1TF U829 ( .A(X_IN[10]), .B(N783), .Y(N278) );
  AOI211X1TF U830 ( .A0(X_IN[10]), .A1(N783), .B0(X_IN[9]), .C0(N761), .Y(N279) );
  INVX2TF U831 ( .A(Y_IN[9]), .Y(N783) );
  AOI211X1TF U832 ( .A0(X_IN[9]), .A1(N761), .B0(N276), .C0(N275), .Y(N280) );
  AOI21X1TF U833 ( .A0(Y_IN[7]), .A1(N489), .B0(N274), .Y(N275) );
  AOI211X1TF U834 ( .A0(N273), .A1(X_IN[7]), .B0(N272), .C0(N271), .Y(N274) );
  NOR2X1TF U835 ( .A(Y_IN[7]), .B(N489), .Y(N272) );
  AOI21X1TF U836 ( .A0(N193), .A1(N464), .B0(N270), .Y(N273) );
  AOI211X1TF U837 ( .A0(N269), .A1(X_IN[5]), .B0(N268), .C0(N267), .Y(N270) );
  NOR2X1TF U838 ( .A(N193), .B(N464), .Y(N268) );
  AOI211X1TF U839 ( .A0(Y_IN[3]), .A1(N443), .B0(N266), .C0(N265), .Y(N269) );
  AOI211X1TF U840 ( .A0(X_IN[4]), .A1(N730), .B0(N85), .C0(N737), .Y(N265) );
  INVX2TF U841 ( .A(Y_IN[3]), .Y(N730) );
  OAI32X1TF U842 ( .A0(N264), .A1(X_IN[2]), .A2(N314), .B0(X_IN[1]), .B1(N264), 
        .Y(N266) );
  OAI211X1TF U843 ( .A0(Y_IN[3]), .A1(N443), .B0(N263), .C0(N316), .Y(N264) );
  INVX2TF U844 ( .A(Y_IN[0]), .Y(N656) );
  INVX2TF U845 ( .A(Y_IN[1]), .Y(N314) );
  AOI22X1TF U846 ( .A0(N85), .A1(N737), .B0(X_IN[2]), .B1(N315), .Y(N263) );
  INVX2TF U847 ( .A(Y_IN[2]), .Y(N737) );
  INVX2TF U848 ( .A(X_IN[4]), .Y(N443) );
  INVX2TF U849 ( .A(X_IN[6]), .Y(N464) );
  INVX2TF U850 ( .A(X_IN[8]), .Y(N489) );
  NOR2X1TF U851 ( .A(Y_IN[9]), .B(N503), .Y(N276) );
  INVX2TF U852 ( .A(X_IN[10]), .Y(N503) );
  INVX2TF U853 ( .A(Y_IN[8]), .Y(N761) );
  INVX2TF U854 ( .A(Y_IN[10]), .Y(N548) );
  NOR2X1TF U855 ( .A(Y_IN[11]), .B(N302), .Y(N282) );
  INVX2TF U856 ( .A(X_IN[12]), .Y(N302) );
  INVX2TF U857 ( .A(N339), .Y(N385) );
  AOI22X1TF U858 ( .A0(N799), .A1(SUM_AB[2]), .B0(SUM_AB[11]), .B1(N138), .Y(
        N816) );
  INVX2TF U859 ( .A(N309), .Y(N628) );
  OAI21X1TF U860 ( .A0(N171), .A1(N105), .B0(N256), .Y(OPER_A[12]) );
  OAI21X1TF U861 ( .A0(N144), .A1(N104), .B0(N246), .Y(OPER_A[3]) );
  OAI21X1TF U862 ( .A0(N151), .A1(N105), .B0(N247), .Y(OPER_A[4]) );
  OAI21X1TF U863 ( .A0(N145), .A1(N105), .B0(N248), .Y(OPER_A[5]) );
  OAI21X1TF U864 ( .A0(N154), .A1(N105), .B0(N249), .Y(OPER_A[6]) );
  OAI21X1TF U865 ( .A0(N143), .A1(N105), .B0(N250), .Y(OPER_A[7]) );
  OAI21X1TF U866 ( .A0(N176), .A1(N105), .B0(N251), .Y(OPER_A[8]) );
  OAI21X1TF U867 ( .A0(N105), .A1(N529), .B0(N252), .Y(OPER_A[9]) );
  OAI21X1TF U868 ( .A0(N105), .A1(N147), .B0(N253), .Y(OPER_A[10]) );
  OAI21X1TF U869 ( .A0(N105), .A1(N155), .B0(N254), .Y(OPER_A[11]) );
  OAI21X1TF U870 ( .A0(N152), .A1(N104), .B0(N245), .Y(OPER_A[2]) );
  INVX2TF U871 ( .A(N559), .Y(N799) );
  NOR2X1TF U872 ( .A(N339), .B(N370), .Y(ALU_IS_DONE) );
  OAI211X1TF U873 ( .A0(N152), .A1(N87), .B0(N223), .C0(N222), .Y(FOUT[0]) );
  AOI31X1TF U874 ( .A0(X_IN[0]), .A1(N119), .A2(N153), .B0(N391), .Y(N392) );
  AOI21X1TF U875 ( .A0(N119), .A1(N473), .B0(N472), .Y(N474) );
  AOI22X1TF U876 ( .A0(N118), .A1(N466), .B0(SUM_AB[8]), .B1(N127), .Y(N468)
         );
  AOI22X1TF U877 ( .A0(N119), .A1(\INTADD_0_SUM[0] ), .B0(SUM_AB[1]), .B1(N130), .Y(N403) );
  AOI22X1TF U878 ( .A0(N119), .A1(\INTADD_0_SUM[3] ), .B0(SUM_AB[4]), .B1(N130), .Y(N432) );
  AOI22X1TF U879 ( .A0(N119), .A1(\INTADD_0_SUM[5] ), .B0(N799), .B1(
        SUM_AB[10]), .Y(N449) );
  AOI31X1TF U880 ( .A0(N118), .A1(N147), .A2(N495), .B0(N490), .Y(N491) );
  AOI22X1TF U881 ( .A0(N119), .A1(\INTADD_0_SUM[1] ), .B0(SUM_AB[2]), .B1(N130), .Y(N413) );
  AOI21X1TF U882 ( .A0(N119), .A1(N357), .B0(N514), .Y(N358) );
  AOI31X1TF U883 ( .A0(N119), .A1(N155), .A2(N511), .B0(N509), .Y(N513) );
  AOI22X1TF U884 ( .A0(N119), .A1(\INTADD_0_SUM[6] ), .B0(SUM_AB[7]), .B1(N130), .Y(N462) );
  AOI22X1TF U885 ( .A0(N118), .A1(\INTADD_0_SUM[4] ), .B0(SUM_AB[5]), .B1(N127), .Y(N439) );
  AOI22X1TF U886 ( .A0(N119), .A1(\INTADD_0_SUM[2] ), .B0(SUM_AB[3]), .B1(N130), .Y(N423) );
  NOR2X1TF U887 ( .A(ALU_TYPE[2]), .B(ALU_TYPE[0]), .Y(N197) );
  NAND3X1TF U888 ( .A(N905), .B(N215), .C(N214), .Y(N674) );
  NAND4BX1TF U889 ( .AN(N838), .B(N210), .C(N839), .D(N209), .Y(N680) );
  AOI2BB2X1TF U890 ( .B0(N107), .B1(C152_DATA4_2), .A0N(N156), .A1N(N929), .Y(
        N209) );
  OAI2BB1X1TF U891 ( .A0N(N107), .A1N(C152_DATA4_10), .B0(N216), .Y(N672) );
  NAND3X1TF U892 ( .A(N866), .B(N867), .C(N212), .Y(N677) );
  OAI2BB2XLTF U893 ( .B0(OFFSET[0]), .B1(N202), .A0N(Y_IN[2]), .A1N(N125), .Y(
        C2_Z_2) );
  AOI2BB2X1TF U894 ( .B0(N220), .B1(DIVISION_REMA[0]), .A0N(N172), .A1N(N81), 
        .Y(N223) );
  OAI222X1TF U895 ( .A0(N97), .A1(N529), .B0(N81), .B1(N163), .C0(N155), .C1(
        N87), .Y(FOUT[9]) );
  NAND2X1TF U896 ( .A(N149), .B(N165), .Y(N370) );
  NAND3X1TF U897 ( .A(STEP[2]), .B(STEP[3]), .C(N643), .Y(N940) );
  NAND3X1TF U898 ( .A(N546), .B(N387), .C(N635), .Y(N648) );
  NOR4XLTF U899 ( .A(N762), .B(N618), .C(N801), .D(N648), .Y(N262) );
  AOI222XLTF U900 ( .A0(STEP[2]), .A1(N150), .B0(N121), .B1(N165), .C0(N142), 
        .C1(N122), .Y(N260) );
  NAND3X1TF U901 ( .A(N262), .B(N361), .C(N634), .Y(N620) );
  AOI2BB1X1TF U902 ( .A0N(X_IN[5]), .A1N(N269), .B0(Y_IN[4]), .Y(N267) );
  AOI2BB1X1TF U903 ( .A0N(X_IN[7]), .A1N(N273), .B0(Y_IN[6]), .Y(N271) );
  NAND2X1TF U904 ( .A(MODE_TYPE[0]), .B(N312), .Y(N763) );
  AO22X1TF U905 ( .A0(X_IN[4]), .A1(N737), .B0(N85), .B1(N315), .Y(N284) );
  NAND2X1TF U906 ( .A(N101), .B(N730), .Y(N286) );
  AOI2BB1X1TF U907 ( .A0N(N290), .A1N(X_IN[6]), .B0(Y_IN[4]), .Y(N288) );
  AOI2BB1X1TF U908 ( .A0N(N294), .A1N(X_IN[8]), .B0(Y_IN[6]), .Y(N292) );
  NAND2X1TF U909 ( .A(N157), .B(N181), .Y(N617) );
  NAND4BX1TF U910 ( .AN(N383), .B(N313), .C(N803), .D(N361), .Y(N725) );
  NAND2X1TF U911 ( .A(N833), .B(N156), .Y(N841) );
  NAND2X1TF U912 ( .A(N852), .B(N177), .Y(N861) );
  NOR2BX1TF U913 ( .AN(N887), .B(OPER_B[7]), .Y(N895) );
  NAND2X1TF U914 ( .A(N895), .B(N160), .Y(N908) );
  NAND2X1TF U915 ( .A(N923), .B(N161), .Y(N936) );
  NAND2X1TF U916 ( .A(N907), .B(N74), .Y(N958) );
  NAND2X1TF U917 ( .A(N566), .B(N958), .Y(N939) );
  NAND2X1TF U918 ( .A(N967), .B(N378), .Y(N574) );
  NAND3X1TF U919 ( .A(N92), .B(N91), .C(N90), .Y(N592) );
  NOR2BX1TF U920 ( .AN(N574), .B(N606), .Y(N571) );
  NAND2X1TF U921 ( .A(PRE_WORK), .B(N351), .Y(N953) );
  NAND2X1TF U922 ( .A(N606), .B(N823), .Y(N344) );
  NAND2X1TF U923 ( .A(N219), .B(N959), .Y(N363) );
  NAND3X1TF U924 ( .A(SIGN_Y), .B(N74), .C(N906), .Y(N824) );
  NAND2X1TF U925 ( .A(N856), .B(N849), .Y(N862) );
  NAND2X1TF U926 ( .A(N875), .B(N876), .Y(N891) );
  NAND2X1TF U927 ( .A(N897), .B(N898), .Y(N909) );
  NAND2X1TF U928 ( .A(N915), .B(N917), .Y(N933) );
  NAND3X1TF U929 ( .A(N606), .B(N603), .C(N162), .Y(N601) );
  NAND2X1TF U930 ( .A(N416), .B(N415), .Y(N424) );
  NAND2X1TF U931 ( .A(N434), .B(N433), .Y(N444) );
  NAND2X1TF U932 ( .A(N454), .B(N453), .Y(N463) );
  NAND2X1TF U933 ( .A(N500), .B(N499), .Y(N1014) );
  AOI222XLTF U934 ( .A0(XTEMP[11]), .A1(X_IN[11]), .B0(XTEMP[11]), .B1(N498), 
        .C0(X_IN[11]), .C1(N498), .Y(N352) );
  XOR2X1TF U935 ( .A(X_IN[12]), .B(N352), .Y(N357) );
  NAND3X1TF U936 ( .A(N567), .B(POST_WORK), .C(N603), .Y(N373) );
  NAND3BX1TF U937 ( .AN(N363), .B(N949), .C(N967), .Y(N599) );
  NAND3X1TF U938 ( .A(N610), .B(N364), .C(N599), .Y(N943) );
  NAND2X1TF U939 ( .A(N112), .B(N395), .Y(N382) );
  NAND3X1TF U940 ( .A(N385), .B(N122), .C(DP_OP_333_124_4748_N57), .Y(N639) );
  NOR2BX1TF U941 ( .AN(N635), .B(N944), .Y(N543) );
  NAND3X1TF U942 ( .A(N543), .B(N377), .C(N376), .Y(N381) );
  NAND4X1TF U943 ( .A(N428), .B(N427), .C(N426), .D(N425), .Y(N429) );
  NAND4X1TF U944 ( .A(N439), .B(N438), .C(N437), .D(N436), .Y(N440) );
  NAND4X1TF U945 ( .A(N449), .B(N448), .C(N447), .D(N446), .Y(N450) );
  OAI2BB1X1TF U946 ( .A0N(DIVISION_HEAD[10]), .A1N(N472), .B0(N452), .Y(N713)
         );
  AOI2BB2X1TF U947 ( .B0(X_IN[9]), .B1(N479), .A0N(N479), .A1N(X_IN[9]), .Y(
        N484) );
  NAND3X1TF U948 ( .A(N118), .B(N529), .C(N484), .Y(N480) );
  AOI2BB1X1TF U949 ( .A0N(N510), .A1N(N484), .B0(N514), .Y(N485) );
  AOI2BB2X1TF U950 ( .B0(N488), .B1(N503), .A0N(N503), .A1N(N488), .Y(N495) );
  AOI2BB1X1TF U951 ( .A0N(N510), .A1N(N495), .B0(N514), .Y(N496) );
  AOI2BB2X1TF U952 ( .B0(N79), .B1(N498), .A0N(N498), .A1N(N79), .Y(N511) );
  OAI2BB2XLTF U953 ( .B0(N503), .B1(N609), .A0N(XTEMP[12]), .A1N(N88), .Y(N504) );
  AOI2BB1X1TF U954 ( .A0N(N510), .A1N(N511), .B0(N514), .Y(N512) );
  AOI2BB1X1TF U955 ( .A0N(DIVISION_REMA[2]), .A1N(N518), .B0(DIVISION_HEAD[6]), 
        .Y(N516) );
  OA21XLTF U956 ( .A0(N151), .A1(DIVISION_REMA[4]), .B0(N520), .Y(N522) );
  OA21XLTF U957 ( .A0(N154), .A1(DIVISION_REMA[6]), .B0(N524), .Y(N526) );
  OA21XLTF U958 ( .A0(XTEMP[12]), .A1(N536), .B0(N148), .Y(N535) );
  NAND4X1TF U959 ( .A(N546), .B(N545), .C(N639), .D(N544), .Y(N557) );
  NAND3X1TF U960 ( .A(N552), .B(N551), .C(N550), .Y(N553) );
  NAND3X1TF U961 ( .A(N756), .B(N560), .C(N559), .Y(N561) );
  NAND3X1TF U962 ( .A(N567), .B(N603), .C(N822), .Y(N573) );
  NAND4X1TF U963 ( .A(N569), .B(N568), .C(N640), .D(N573), .Y(N570) );
  NAND2X1TF U964 ( .A(N180), .B(N158), .Y(N591) );
  NOR4XLTF U965 ( .A(\RSHT_BITS[3] ), .B(N90), .C(N615), .D(N591), .Y(N572) );
  NAND2X1TF U966 ( .A(N580), .B(N590), .Y(N587) );
  NAND2X1TF U967 ( .A(N92), .B(N91), .Y(N589) );
  AOI2BB2X1TF U968 ( .B0(N597), .B1(N158), .A0N(N591), .A1N(N593), .Y(N585) );
  NAND4X1TF U969 ( .A(N94), .B(N635), .C(N634), .D(N633), .Y(N636) );
  NAND4X1TF U970 ( .A(N641), .B(N640), .C(N639), .D(N644), .Y(N697) );
  NAND3X1TF U971 ( .A(N756), .B(N652), .C(N651), .Y(N653) );
  AO22X1TF U972 ( .A0(DIVISION_REMA[4]), .A1(N735), .B0(N193), .B1(N790), .Y(
        N743) );
  AOI2BB1X1TF U973 ( .A0N(X_IN[1]), .A1N(N764), .B0(N763), .Y(N767) );
  NAND4X1TF U974 ( .A(N794), .B(N793), .C(N792), .D(N791), .Y(N795) );
  OAI221XLTF U975 ( .A0(\INDEX[2] ), .A1(N90), .B0(N124), .B1(\RSHT_BITS[3] ), 
        .C0(N817), .Y(N818) );
  OAI221XLTF U976 ( .A0(N129), .A1(N180), .B0(N157), .B1(N92), .C0(N819), .Y(
        N830) );
  NAND2X1TF U977 ( .A(N904), .B(N870), .Y(N865) );
  NAND2BX1TF U978 ( .AN(N820), .B(N865), .Y(N886) );
  NAND2X1TF U979 ( .A(N829), .B(N967), .Y(N871) );
  NAND3X1TF U980 ( .A(SIGN_Y), .B(N74), .C(N221), .Y(N837) );
  OAI2BB1X1TF U981 ( .A0N(N960), .A1N(N830), .B0(N829), .Y(N920) );
  NAND3X1TF U982 ( .A(N74), .B(N178), .C(N56), .Y(N975) );
  NAND4X1TF U983 ( .A(N221), .B(N178), .C(N56), .D(N965), .Y(N839) );
  NAND2X1TF U984 ( .A(N904), .B(N920), .Y(N938) );
  NAND3BX1TF U985 ( .AN(OPER_A[7]), .B(N931), .C(N891), .Y(N892) );
  NAND2X1TF U986 ( .A(N941), .B(N946), .Y(N947) );
  NAND2X1TF U987 ( .A(N979), .B(N978), .Y(N668) );
  NAND2X1TF U988 ( .A(N982), .B(N981), .Y(N667) );
  NAND2X1TF U989 ( .A(SUM_AB[3]), .B(N83), .Y(N983) );
  NAND2X1TF U990 ( .A(N988), .B(N987), .Y(N665) );
  NAND2X1TF U991 ( .A(SUM_AB[5]), .B(N83), .Y(N989) );
  NAND2X1TF U992 ( .A(N994), .B(N993), .Y(N663) );
  NAND2X1TF U993 ( .A(SUM_AB[7]), .B(N83), .Y(N995) );
  NAND2X1TF U994 ( .A(N1000), .B(N999), .Y(N661) );
  NAND2X1TF U995 ( .A(SUM_AB[9]), .B(N83), .Y(N1001) );
  NAND2X1TF U996 ( .A(N1006), .B(N1005), .Y(N659) );
  NAND2X1TF U997 ( .A(SUM_AB[11]), .B(N83), .Y(N1007) );
endmodule


module SERIAL_CPU_8BIT_VG ( CLK, ENABLE, RST_N, START, I_DATAIN, D_DATAIN, 
        IS_I_ADDR, NXT, I_ADDR, D_ADDR, D_WE, D_DATAOUT, IO_STATUS, IO_CONTROL, 
        IO_DATAINA, IO_DATAINB, IO_DATAOUTA, IO_DATAOUTB, IO_OFFSET );
  input [7:0] I_DATAIN;
  input [7:0] D_DATAIN;
  output [1:0] NXT;
  output [8:0] I_ADDR;
  output [8:0] D_ADDR;
  output [7:0] D_DATAOUT;
  input [15:0] IO_STATUS;
  output [15:0] IO_CONTROL;
  input [15:0] IO_DATAINA;
  input [15:0] IO_DATAINB;
  output [15:0] IO_DATAOUTA;
  output [15:0] IO_DATAOUTB;
  output [15:0] IO_OFFSET;
  input CLK, ENABLE, RST_N, START;
  output IS_I_ADDR, D_WE;
  wire   \OPER1_R1[2] , N110, N166, N167, N168, CF_BUF, N470, N471, N472, N473,
         N474, N475, N476, N477, N478, N479, N480, N481, N482, N483, N484,
         N485, N486, N504, N505, N506, N507, N508, N509, N510, N511, N512,
         N513, N514, N515, N516, N517, N518, N519, N588, N589, ZF, CF, N616,
         N400, N401, N402, N403, N404, N405, N406, N408, N409, N411, N412,
         N413, N414, N415, N416, N418, N420, N421, N423, N424, N433, N434,
         N435, N436, N437, N438, N439, N440, N441, N442, N443, N444, N445,
         N447, N448, N449, N451, N452, N453, N455, N456, N457, N459, N460,
         N461, N462, N464, N465, N466, N468, N469, N4700, N4720, N4730, N4740,
         N4750, N4770, N4780, N4790, N4800, N4820, N4830, N4840, N4860, N487,
         N488, N489, N491, N492, N493, N495, N496, N497, N498, N500, N501,
         N502, N503, N5050, N5060, N5070, N5080, N5100, N5110, N5130, N5140,
         N5180, N520, N521, N522, N523, N524, N525, N526, N527, N528, N529,
         N530, N531, N532, N533, N534, N535, N554, N569, N571, N572, N595,
         N596, N597, N598, N599, N600, N601, N602, N603, N604, N605, N606,
         N607, N608, N609, N610, N613, N614, N615, N6160, N617, N618, N619,
         N620, N621, N622, N623, N624, N625, N626, N627, N628, N629, N630,
         N631, N632, N633, N634, N635, N636, N637, N638, N639, N640, N641,
         N642, N643, N644, N645, N646, N647, N648, N649, N650, N651, N652,
         N653, N654, N655, N656, N657, N658, N659, N660, N661, N662, N663,
         N664, N665, N666, N667, N668, N669, N670, N671, N672, N673, N674,
         N675, N676, N677, N678, N679, N680, N681, N682, N683, N684, N685,
         N686, N687, N688, N689, N690, N691, N692, N804, N808, N809, N810,
         N811, N812, N859, N860, N922, N923, N924, N925, N926, N927, N928,
         N929, N930, N931, N932, N933, N934, N935, N936, N937, N938, N939,
         N940, N941, N942, N943, N944, N945, N946, N947, N948, N949, N950,
         N951, N952, N953, N954, N955, N956, N957, N958, N959, N960, N961,
         N962, N963, N964, N965, N966, N967, N968, N969, N970, N971, N972,
         N973, N974, N975, N976, N977, N978, N979, N980, N981, N982, N983,
         N984, N985, N986, N987, N988, N989, N990, N991, N992, N993, N994,
         N995, N996, N997, N998, N999, N1000, N1001, N1002, SUB_X_285_4_N16,
         SUB_X_285_4_N15, SUB_X_285_4_N14, SUB_X_285_4_N13, SUB_X_285_4_N12,
         SUB_X_285_4_N11, SUB_X_285_4_N10, SUB_X_285_4_N9, SUB_X_285_4_N8,
         SUB_X_285_4_N7, SUB_X_285_4_N6, SUB_X_285_4_N5, SUB_X_285_4_N4,
         SUB_X_285_4_N3, SUB_X_285_4_N2, SUB_X_285_4_N1, ADD_X_285_3_N16,
         ADD_X_285_3_N15, ADD_X_285_3_N14, ADD_X_285_3_N13, ADD_X_285_3_N12,
         ADD_X_285_3_N11, ADD_X_285_3_N10, ADD_X_285_3_N9, ADD_X_285_3_N8,
         ADD_X_285_3_N7, ADD_X_285_3_N6, ADD_X_285_3_N5, ADD_X_285_3_N4,
         ADD_X_285_3_N3, ADD_X_285_3_N2, N1, N2, N3, N4, N5, N6, N7, N8, N9,
         N10, N11, N12, N13, N14, N15, N16, N17, N18, N19, N20, N21, N22, N23,
         N24, N25, N26, N35, N121, N122, N123, N124, N125, N126, N127, N128,
         N129, N130, N131, N132, N133, N134, N135, N136, N137, N138, N139,
         N140, N141, N142, N143, N144, N145, N146, N147, N148, N149, N150,
         N151, N152, N153, N154, N155, N156, N157, N158, N159, N160, N161,
         N162, N163, N164, N165, N1660, N1670, N1680, N169, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200,
         N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211,
         N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222,
         N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233,
         N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244,
         N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255,
         N256, N257, N258, N259, N260, N261, N262, N263, N264, N265, N266,
         N267, N268, N269, N270, N271, N272, N273, N274, N275, N276, N277,
         N278, N279, N280, N281, N282, N283, N284, N285, N286, N287, N288,
         N289, N290, N291, N292, N293, N294, N295, N296, N297, N298, N299,
         N300, N301, N302, N303, N304, N305, N306, N307, N308, N309, N310,
         N311, N312, N313, N314, N315, N316, N317, N318, N319, N320, N321,
         N322, N323, N324, N325, N326, N327, N328, N329, N330, N331, N332,
         N333, N334, N335, N336, N337, N338, N339, N340, N341, N342, N343,
         N344, N345, N346, N347, N348, N349, N350, N351, N352, N353, N354,
         N355, N356, N357, N358, N359, N360, N361, N362, N363, N364, N365,
         N366, N367, N368, N369, N370, N371, N372, N373, N374, N375, N376,
         N377, N378, N379, N380, N381, N382, N383, N384, N385, N386, N387,
         N388, N389, N390, N391, N392, N393, N394, N395, N396, N397, N398,
         N399, N407, N410, N417, N419, N422, N425, N426, N427, N428, N429,
         N430, N431, N432, N446, N450, N454, N458, N463, N467, N4710, N4760,
         N4810, N4850, N490, N494, N499, N5040, N5090, N5120, N5150, N5160,
         N5170, N5190, N536, N537, N538, N539, N540, N541, N542, N543, N544,
         N545, N546, N547, N548, N549, N550, N551, N552, N553, N555, N556,
         N557, N558, N559, N560, N561, N562, N563, N564, N565, N566, N567,
         N568, N570, N573, N574, N575, N576, N577, N578, N579, N580, N581,
         N582, N583, N584, N585, N586, N587, N5880, N5890, N590, N591, N592,
         N593, N594, N611, N612, N693, N694, N695, N696, N697, N698, N699,
         N700, N701, N702, N703, N704, N705, N706, N707, N708, N709, N710,
         N711, N712, N713, N714, N715, N716, N717, N718, N719, N720, N721,
         N722, N723, N724, N725, N726, N727, N728, N729, N730, N731, N732,
         N733, N734, N735, N736, N737, N738, N739, N740, N741, N742, N743,
         N744, N745, N746, N747, N748, N749, N750, N751, N752, N753, N754,
         N755, N756, N757, N758, N759, N760, N761, N762, N763, N764, N765,
         N766, N767, N768, N769, N770, N771, N772, N773, N774, N775, N776,
         N777, N778, N779, N780, N781, N782, N783, N784, N785, N786, N787,
         N788, N789, N790, N791, N792, N793, N794, N795, N796, N797, N798,
         N799, N800, N801, N802, N803, N805, N806, N807, N813, N814, N815,
         N816, N817, N818, N819, N820, N821, N822, N823, N824, N825, N826,
         N827, N828, N829, N830, N831, N832, N833, N834, N835, N836, N837,
         N838, N839, N840, N841, N842, N843, N844, N845, N846, N847, N848,
         N849, N850, N851, N852, N853, N854, N855, N856, N857, N858, N861,
         N862, N863, N864, N865, N866, N867, N868, N869, N870, N871, N872,
         N873, N874, N875, N876, N877, N878, N879, N880, N881, N882, N883,
         N884, N885, N886, N887, N888, N889, N890, N891, N892, N893, N894,
         N895, N896, N897, N898, N899, N900, N901, N902, N903, N904, N905,
         N906, N907, N908, N909, N910, N911, N912, N913, N914, N915, N916,
         N917, N918, N919, N920, N921, N1003, N1004, N1005, N1006, N1007,
         N1008, N1009, N1010, N1011, N1012, N1013, N1014, N1015, N1016, N1017,
         N1018, N1019, N1020, N1021, N1022, N1023, N1024, N1025, N1026, N1027,
         N1028, N1029, N1030, N1031, N1032, N1033, N1034, N1035, N1036, N1037,
         N1038, N1039, N1040, N1041, N1042, N1043, N1044, N1045, N1046, N1047,
         N1048, N1049, N1050, N1051, N1052, N1053, N1054, N1055, N1056, N1057,
         N1058, N1059, N1060, N1061, N1062, N1063, N1064, N1065, N1066, N1067,
         N1068, N1069, N1070, N1071, N1072, N1073, N1074, N1075, N1076, N1077,
         N1078, N1079, N1080, N1081, N1082, N1083, N1084, N1085, N1086, N1087,
         N1088, N1089, N1090, N1091, N1092, N1093, N1094, N1095, N1096, N1097,
         N1098, N1099, N11000, N1101, N1102, N1103, N1104, N1105, N1106, N1107,
         N1108, N1109, N1110, N1111, N1112, N1113, N1114, N1115, N1116, N1117,
         N1118, N1119, N1120, N1121, N1122, N1123, N1124, N1125, N1126, N1127,
         N1128, N1129, N1130, N1131, N1132, N1133, N1134, N1135, N1136, N1137,
         N1138, N1139, N1140, N1141, N1142, N1143, N1144, N1145, N1146, N1147,
         N1148, N1149, N1150, N1151, N1152, N1153, N1154, N1155, N1156, N1157,
         N1158, N1159, N1160, N1161, N1162, N1163, N1164, N1165, N1166, N1167,
         N1168, N1169, N1170, N1171, N1172, N1173, N1174, N1175, N1176, N1177,
         N1178, N1179, N1180, N1181, N1182, N1183, N1184, N1185, N1186, N1187,
         N1188, N1189, N1190, N1191, N1192, N1193;
  wire   [4:2] CODE_TYPE;
  wire   [2:0] OPER3_R3;
  wire   [3:0] STATE;
  wire   [3:0] NEXT_STATE;
  wire   [15:0] REG_A;
  wire   [15:0] REG_B;
  wire   [12:8] REG_C;

  DFFRX4TF \reg_A_reg[0]  ( .D(N497), .CK(CLK), .RN(RST_N), .Q(REG_A[0]), .QN(
        N187) );
  DFFRX4TF \reg_B_reg[1]  ( .D(N487), .CK(CLK), .RN(RST_N), .Q(REG_B[1]), .QN(
        N200) );
  DFFRX2TF \id_ir_reg[11]  ( .D(N532), .CK(CLK), .RN(RST_N), .Q(N186), .QN(
        N569) );
  DFFRX2TF \gr_reg[3][12]  ( .D(N932), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTB[12]), .QN(N632) );
  DFFRX2TF \gr_reg[1][5]  ( .D(N987), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[5]), 
        .QN(N671) );
  DFFRX2TF \gr_reg[3][4]  ( .D(N972), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[4]), 
        .QN(N640) );
  DFFRX2TF \gr_reg[3][6]  ( .D(N970), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[6]), 
        .QN(N638) );
  DFFRX2TF \gr_reg[3][5]  ( .D(N971), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[5]), 
        .QN(N639) );
  DFFRX2TF \gr_reg[1][4]  ( .D(N988), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[4]), 
        .QN(N672) );
  DFFRX2TF \gr_reg[3][11]  ( .D(N933), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTB[11]), .QN(N633) );
  DFFRX2TF \gr_reg[3][0]  ( .D(N976), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[0]), 
        .QN(N644) );
  DFFRX2TF \gr_reg[3][15]  ( .D(N929), .CK(CLK), .RN(RST_N), .Q(N216), .QN(
        N629) );
  DFFRX2TF \gr_reg[3][1]  ( .D(N975), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[1]), 
        .QN(N643) );
  DFFRX2TF \gr_reg[3][14]  ( .D(N930), .CK(CLK), .RN(RST_N), .Q(N215), .QN(
        N630) );
  DFFRX2TF \gr_reg[3][10]  ( .D(N934), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTB[10]), .QN(N634) );
  DFFRX2TF \gr_reg[3][9]  ( .D(N935), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[9]), 
        .QN(N635) );
  DFFRX2TF \gr_reg[3][13]  ( .D(N931), .CK(CLK), .RN(RST_N), .Q(N214), .QN(
        N631) );
  DFFRX2TF \gr_reg[3][2]  ( .D(N974), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[2]), 
        .QN(N642) );
  DFFRX2TF \gr_reg[3][8]  ( .D(N936), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[8]), 
        .QN(N636) );
  DFFRX2TF zf_reg ( .D(N434), .CK(CLK), .RN(RST_N), .Q(ZF), .QN(N213) );
  DFFSX2TF \pc_reg[6]  ( .D(N804), .CK(CLK), .SN(RST_N), .Q(N212), .QN(
        I_ADDR[7]) );
  DFFRX2TF \id_ir_reg[8]  ( .D(N535), .CK(CLK), .RN(RST_N), .Q(N210), .QN(N572) );
  DFFSX2TF \pc_reg[4]  ( .D(N809), .CK(CLK), .SN(RST_N), .Q(N209), .QN(
        I_ADDR[5]) );
  DFFSX2TF \pc_reg[1]  ( .D(N812), .CK(CLK), .SN(RST_N), .Q(N208), .QN(
        I_ADDR[2]) );
  DFFRX2TF \reg_A_reg[6]  ( .D(N448), .CK(CLK), .RN(RST_N), .Q(REG_A[6]), .QN(
        N207) );
  DFFRX2TF \reg_A_reg[8]  ( .D(N456), .CK(CLK), .RN(RST_N), .Q(REG_A[8]), .QN(
        N206) );
  DFFRX2TF \reg_A_reg[4]  ( .D(N452), .CK(CLK), .RN(RST_N), .Q(REG_A[4]), .QN(
        N202) );
  DFFRX2TF \gr_reg[1][6]  ( .D(N986), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[6]), 
        .QN(N670) );
  DFFRX2TF \gr_reg[3][7]  ( .D(N969), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[7]), 
        .QN(N637) );
  DFFRX2TF \id_ir_reg[4]  ( .D(N523), .CK(CLK), .RN(RST_N), .Q(N199), .QN(N401) );
  DFFRX2TF \id_ir_reg[0]  ( .D(N527), .CK(CLK), .RN(RST_N), .Q(OPER3_R3[0]), 
        .QN(N198) );
  DFFRX2TF \id_ir_reg[10]  ( .D(N533), .CK(CLK), .RN(RST_N), .Q(\OPER1_R1[2] ), 
        .QN(N197) );
  DFFSX2TF \pc_reg[0]  ( .D(N860), .CK(CLK), .SN(RST_N), .Q(N196), .QN(
        I_ADDR[1]) );
  DFFRX2TF \state_reg[3]  ( .D(NEXT_STATE[3]), .CK(CLK), .RN(RST_N), .Q(
        STATE[3]), .QN(N195) );
  DFFRX2TF \reg_A_reg[11]  ( .D(N5070), .CK(CLK), .RN(RST_N), .Q(REG_A[11]), 
        .QN(N194) );
  DFFRX2TF \reg_A_reg[15]  ( .D(N492), .CK(CLK), .RN(RST_N), .Q(REG_A[15]), 
        .QN(N192) );
  DFFRX2TF \id_ir_reg[14]  ( .D(N529), .CK(CLK), .RN(RST_N), .Q(CODE_TYPE[3]), 
        .QN(N191) );
  DFFRX2TF \reg_A_reg[12]  ( .D(N502), .CK(CLK), .RN(RST_N), .Q(REG_A[12]), 
        .QN(N190) );
  DFFRX2TF \reg_A_reg[7]  ( .D(N5110), .CK(CLK), .RN(RST_N), .Q(REG_A[7]), 
        .QN(N189) );
  DFFRX2TF \reg_A_reg[10]  ( .D(N4740), .CK(CLK), .RN(RST_N), .Q(REG_A[10]), 
        .QN(N188) );
  DFFRX2TF \id_ir_reg[1]  ( .D(N526), .CK(CLK), .RN(RST_N), .Q(OPER3_R3[1]), 
        .QN(N185) );
  DFFSX2TF \pc_reg[2]  ( .D(N811), .CK(CLK), .SN(RST_N), .Q(N184), .QN(
        I_ADDR[3]) );
  DFFRX2TF \state_reg[1]  ( .D(NEXT_STATE[1]), .CK(CLK), .RN(RST_N), .Q(
        STATE[1]), .QN(N183) );
  DFFRX2TF \id_ir_reg[15]  ( .D(N528), .CK(CLK), .RN(RST_N), .Q(CODE_TYPE[4]), 
        .QN(N182) );
  DFFRX2TF \id_ir_reg[13]  ( .D(N530), .CK(CLK), .RN(RST_N), .Q(CODE_TYPE[2]), 
        .QN(N181) );
  DFFRX2TF \reg_B_reg[3]  ( .D(N4780), .CK(CLK), .RN(RST_N), .Q(REG_B[3]), 
        .QN(N204) );
  DFFRX2TF \id_ir_reg[2]  ( .D(N525), .CK(CLK), .RN(RST_N), .Q(OPER3_R3[2]), 
        .QN(N180) );
  DFFRX2TF \state_reg[2]  ( .D(NEXT_STATE[2]), .CK(CLK), .RN(RST_N), .Q(N179), 
        .QN(N554) );
  DFFRX2TF \reg_A_reg[13]  ( .D(N465), .CK(CLK), .RN(RST_N), .Q(REG_A[13]), 
        .QN(N178) );
  DFFRX2TF \reg_A_reg[9]  ( .D(N469), .CK(CLK), .RN(RST_N), .Q(REG_A[9]), .QN(
        N176) );
  TLATXLTF cf_buf_reg ( .G(N588), .D(N589), .Q(CF_BUF) );
  TLATXLTF \nxt_reg[0]  ( .G(N166), .D(N167), .Q(NXT[0]) );
  TLATXLTF \nxt_reg[1]  ( .G(N166), .D(N168), .Q(NXT[1]) );
  DFFRX2TF \gr_reg[4][9]  ( .D(N927), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[9]), 
        .QN(N619) );
  DFFRX2TF \gr_reg[4][7]  ( .D(N961), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[7]), 
        .QN(N621) );
  DFFRX2TF \gr_reg[4][8]  ( .D(N928), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[8]), 
        .QN(N620) );
  DFFRX2TF \gr_reg[4][6]  ( .D(N962), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[6]), 
        .QN(N622) );
  DFFRX2TF \gr_reg[4][5]  ( .D(N963), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[5]), 
        .QN(N623) );
  DFFRX2TF \gr_reg[4][1]  ( .D(N967), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[1]), 
        .QN(N627) );
  DFFRX2TF \gr_reg[4][3]  ( .D(N965), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[3]), 
        .QN(N625) );
  DFFRX2TF \gr_reg[4][2]  ( .D(N966), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[2]), 
        .QN(N626) );
  DFFRX2TF \gr_reg[4][4]  ( .D(N964), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[4]), 
        .QN(N624) );
  DFFRX2TF \gr_reg[4][0]  ( .D(N968), .CK(CLK), .RN(RST_N), .Q(IO_OFFSET[0]), 
        .QN(N628) );
  DFFSX2TF \pc_reg[5]  ( .D(N808), .CK(CLK), .SN(RST_N), .QN(I_ADDR[6]) );
  DFFSX2TF \pc_reg[7]  ( .D(N859), .CK(CLK), .SN(RST_N), .QN(I_ADDR[8]) );
  DFFSX2TF \pc_reg[3]  ( .D(N810), .CK(CLK), .SN(RST_N), .QN(I_ADDR[4]) );
  DFFRX2TF \gr_reg[1][0]  ( .D(N992), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[0]), 
        .QN(N676) );
  DFFRX2TF \gr_reg[1][1]  ( .D(N991), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[1]), 
        .QN(N675) );
  DFFRX2TF \gr_reg[2][11]  ( .D(N941), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTA[11]), .QN(N649) );
  DFFRX2TF \reg_B_reg[14]  ( .D(N437), .CK(CLK), .RN(RST_N), .Q(REG_B[14]), 
        .QN(N415) );
  DFFRX2TF \reg_B_reg[15]  ( .D(N436), .CK(CLK), .RN(RST_N), .Q(REG_B[15]), 
        .QN(N412) );
  DFFRX2TF \gr_reg[2][12]  ( .D(N940), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTA[12]), .QN(N648) );
  DFFRX2TF \gr_reg[2][8]  ( .D(N944), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[8]), 
        .QN(N652) );
  DFFRX2TF \gr_reg[2][10]  ( .D(N942), .CK(CLK), .RN(RST_N), .Q(
        IO_DATAOUTA[10]), .QN(N650) );
  DFFRX2TF \gr_reg[2][9]  ( .D(N943), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[9]), 
        .QN(N651) );
  DFFRX2TF \reg_B_reg[11]  ( .D(N5060), .CK(CLK), .RN(RST_N), .Q(REG_B[11]), 
        .QN(N409) );
  DFFRX2TF \reg_B_reg[12]  ( .D(N501), .CK(CLK), .RN(RST_N), .Q(REG_B[12]), 
        .QN(N411) );
  DFFRX2TF \reg_B_reg[10]  ( .D(N4730), .CK(CLK), .RN(RST_N), .Q(REG_B[10]), 
        .QN(N408) );
  DFFRX2TF \reg_B_reg[13]  ( .D(N439), .CK(CLK), .RN(RST_N), .Q(REG_B[13]), 
        .QN(N413) );
  DFFRX2TF \reg_B_reg[9]  ( .D(N438), .CK(CLK), .RN(RST_N), .Q(REG_B[9]), .QN(
        N418) );
  DFFRX2TF \gr_reg[2][3]  ( .D(N981), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[3]), 
        .QN(N657) );
  DFFRX2TF \gr_reg[2][5]  ( .D(N979), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[5]), 
        .QN(N655) );
  DFFRX2TF \gr_reg[1][2]  ( .D(N990), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[2]), 
        .QN(N674) );
  DFFRX2TF \gr_reg[1][3]  ( .D(N989), .CK(CLK), .RN(RST_N), .Q(IO_CONTROL[3]), 
        .QN(N673) );
  DFFRX2TF \gr_reg[2][1]  ( .D(N983), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[1]), 
        .QN(N659) );
  DFFRX2TF \gr_reg[2][6]  ( .D(N978), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[6]), 
        .QN(N654) );
  DFFRX2TF \gr_reg[2][2]  ( .D(N982), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[2]), 
        .QN(N658) );
  DFFRX2TF \state_reg[0]  ( .D(NEXT_STATE[0]), .CK(CLK), .RN(RST_N), .Q(
        STATE[0]), .QN(N205) );
  DFFRX2TF \gr_reg[2][7]  ( .D(N977), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[7]), 
        .QN(N653) );
  DFFRX2TF \gr_reg[2][4]  ( .D(N980), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[4]), 
        .QN(N656) );
  DFFRX2TF \reg_B_reg[7]  ( .D(N5140), .CK(CLK), .RN(RST_N), .Q(REG_B[7]), 
        .QN(N405) );
  DFFRX2TF \reg_B_reg[5]  ( .D(N443), .CK(CLK), .RN(RST_N), .Q(REG_B[5]), .QN(
        N424) );
  DFFRX2TF \reg_B_reg[6]  ( .D(N442), .CK(CLK), .RN(RST_N), .Q(REG_B[6]), .QN(
        N406) );
  DFFRX2TF \reg_B_reg[8]  ( .D(N440), .CK(CLK), .RN(RST_N), .Q(REG_B[8]), .QN(
        N420) );
  DFFRX2TF \gr_reg[2][0]  ( .D(N984), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTA[0]), 
        .QN(N660) );
  DFFRX2TF \gr_reg[3][3]  ( .D(N973), .CK(CLK), .RN(RST_N), .Q(IO_DATAOUTB[3]), 
        .QN(N641) );
  DFFRX2TF \reg_B_reg[4]  ( .D(N441), .CK(CLK), .RN(RST_N), .Q(REG_B[4]), .QN(
        N423) );
  CMPR32X2TF \sub_x_285_4/U15  ( .A(N201), .B(REG_A[2]), .C(SUB_X_285_4_N15), 
        .CO(SUB_X_285_4_N14), .S(N506) );
  CMPR32X2TF \sub_x_285_4/U10  ( .A(N405), .B(REG_A[7]), .C(SUB_X_285_4_N10), 
        .CO(SUB_X_285_4_N9), .S(N511) );
  CMPR32X2TF \sub_x_285_4/U9  ( .A(N420), .B(REG_A[8]), .C(SUB_X_285_4_N9), 
        .CO(SUB_X_285_4_N8), .S(N512) );
  CMPR32X2TF \sub_x_285_4/U8  ( .A(N418), .B(REG_A[9]), .C(SUB_X_285_4_N8), 
        .CO(SUB_X_285_4_N7), .S(N513) );
  CMPR32X2TF \sub_x_285_4/U7  ( .A(N408), .B(REG_A[10]), .C(SUB_X_285_4_N7), 
        .CO(SUB_X_285_4_N6), .S(N514) );
  CMPR32X2TF \sub_x_285_4/U6  ( .A(N409), .B(REG_A[11]), .C(SUB_X_285_4_N6), 
        .CO(SUB_X_285_4_N5), .S(N515) );
  CMPR32X2TF \sub_x_285_4/U5  ( .A(N411), .B(REG_A[12]), .C(SUB_X_285_4_N5), 
        .CO(SUB_X_285_4_N4), .S(N516) );
  CMPR32X2TF \sub_x_285_4/U4  ( .A(N413), .B(REG_A[13]), .C(SUB_X_285_4_N4), 
        .CO(SUB_X_285_4_N3), .S(N517) );
  CMPR32X2TF \sub_x_285_4/U3  ( .A(N415), .B(REG_A[14]), .C(SUB_X_285_4_N3), 
        .CO(SUB_X_285_4_N2), .S(N518) );
  CMPR32X2TF \add_x_285_3/U5  ( .A(REG_A[12]), .B(REG_B[12]), .C(
        ADD_X_285_3_N5), .CO(ADD_X_285_3_N4), .S(N482) );
  CMPR32X2TF \add_x_285_3/U6  ( .A(REG_A[11]), .B(REG_B[11]), .C(
        ADD_X_285_3_N6), .CO(ADD_X_285_3_N5), .S(N481) );
  CMPR32X2TF \add_x_285_3/U7  ( .A(REG_A[10]), .B(REG_B[10]), .C(
        ADD_X_285_3_N7), .CO(ADD_X_285_3_N6), .S(N480) );
  CMPR32X2TF \add_x_285_3/U3  ( .A(REG_A[14]), .B(REG_B[14]), .C(
        ADD_X_285_3_N3), .CO(ADD_X_285_3_N2), .S(N484) );
  CMPR32X2TF \add_x_285_3/U15  ( .A(REG_A[2]), .B(REG_B[2]), .C(
        ADD_X_285_3_N15), .CO(ADD_X_285_3_N14), .S(N472) );
  CMPR32X2TF \add_x_285_3/U13  ( .A(REG_A[4]), .B(REG_B[4]), .C(
        ADD_X_285_3_N13), .CO(ADD_X_285_3_N12), .S(N474) );
  CMPR32X2TF \add_x_285_3/U12  ( .A(REG_A[5]), .B(REG_B[5]), .C(
        ADD_X_285_3_N12), .CO(ADD_X_285_3_N11), .S(N475) );
  CMPR32X2TF \add_x_285_3/U11  ( .A(REG_A[6]), .B(REG_B[6]), .C(
        ADD_X_285_3_N11), .CO(ADD_X_285_3_N10), .S(N476) );
  CMPR32X2TF \add_x_285_3/U10  ( .A(REG_A[7]), .B(REG_B[7]), .C(
        ADD_X_285_3_N10), .CO(ADD_X_285_3_N9), .S(N477) );
  CMPR32X2TF \add_x_285_3/U9  ( .A(REG_A[8]), .B(REG_B[8]), .C(ADD_X_285_3_N9), 
        .CO(ADD_X_285_3_N8), .S(N478) );
  CMPR32X2TF \add_x_285_3/U8  ( .A(REG_A[9]), .B(REG_B[9]), .C(ADD_X_285_3_N8), 
        .CO(ADD_X_285_3_N7), .S(N479) );
  CMPR32X2TF \add_x_285_3/U4  ( .A(REG_A[13]), .B(REG_B[13]), .C(
        ADD_X_285_3_N4), .CO(ADD_X_285_3_N3), .S(N483) );
  DFFNSRX2TF lowest_bit_reg ( .D(N1002), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        I_ADDR[0]), .QN(N193) );
  DFFNSRXLTF is_i_addr_reg ( .D(N110), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        IS_I_ADDR) );
  DFFNSRXLTF dw_reg ( .D(N616), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(D_WE) );
  DFFNSRXLTF \reg_C_reg[12]  ( .D(N5050), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        REG_C[12]) );
  DFFNSRXLTF \reg_C_reg[11]  ( .D(N5100), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        REG_C[11]) );
  DFFNSRXLTF \reg_C_reg[9]  ( .D(N4720), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        REG_C[9]) );
  DFFNSRXLTF \reg_C_reg[8]  ( .D(N459), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        REG_C[8]) );
  DFFNSRXLTF \reg_C_reg[10]  ( .D(N4770), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        REG_C[10]) );
  DFFNSRXLTF \reg_C_reg[13]  ( .D(N468), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N421) );
  DFFNSRXLTF \reg_C_reg[15]  ( .D(N495), .CKN(CLK), .SN(1'b1), .RN(1'b1), .QN(
        N414) );
  DFFNSRXLTF \reg_C_reg[14]  ( .D(N4860), .CKN(CLK), .SN(1'b1), .RN(1'b1), 
        .QN(N416) );
  DFFRX2TF \reg_A_reg[1]  ( .D(N488), .CK(CLK), .RN(RST_N), .Q(REG_A[1]), .QN(
        N1112) );
  DFFRX2TF \reg_A_reg[2]  ( .D(N461), .CK(CLK), .RN(RST_N), .Q(REG_A[2]), .QN(
        N177) );
  DFFRX1TF \smdr_reg[15]  ( .D(N493), .CK(CLK), .RN(RST_N), .QN(N595) );
  DFFRX1TF \smdr_reg[10]  ( .D(N4750), .CK(CLK), .RN(RST_N), .QN(N600) );
  DFFRX1TF \smdr_reg[8]  ( .D(N457), .CK(CLK), .RN(RST_N), .QN(N602) );
  DFFRX1TF \smdr_reg[4]  ( .D(N453), .CK(CLK), .RN(RST_N), .QN(N606) );
  DFFRX1TF \smdr_reg[3]  ( .D(N4800), .CK(CLK), .RN(RST_N), .QN(N607) );
  DFFRX1TF \smdr_reg[0]  ( .D(N498), .CK(CLK), .RN(RST_N), .QN(N610) );
  DFFRX1TF \smdr_reg[1]  ( .D(N489), .CK(CLK), .RN(RST_N), .QN(N609) );
  DFFRX1TF \smdr_reg[14]  ( .D(N4840), .CK(CLK), .RN(RST_N), .QN(N596) );
  DFFRX1TF \smdr_reg[13]  ( .D(N466), .CK(CLK), .RN(RST_N), .QN(N597) );
  DFFRX1TF \smdr_reg[12]  ( .D(N503), .CK(CLK), .RN(RST_N), .QN(N598) );
  DFFRX1TF \smdr_reg[11]  ( .D(N5080), .CK(CLK), .RN(RST_N), .QN(N599) );
  DFFRX1TF \smdr_reg[9]  ( .D(N4700), .CK(CLK), .RN(RST_N), .QN(N601) );
  DFFRX1TF \smdr_reg[7]  ( .D(N433), .CK(CLK), .RN(RST_N), .QN(N603) );
  DFFRX1TF \smdr_reg[6]  ( .D(N449), .CK(CLK), .RN(RST_N), .QN(N604) );
  DFFRX1TF \smdr_reg[5]  ( .D(N445), .CK(CLK), .RN(RST_N), .QN(N605) );
  DFFRX1TF \smdr_reg[2]  ( .D(N462), .CK(CLK), .RN(RST_N), .QN(N608) );
  DFFRX1TF nf_reg ( .D(N435), .CK(CLK), .RN(RST_N), .QN(N211) );
  DFFRX1TF \id_ir_reg[7]  ( .D(N520), .CK(CLK), .RN(RST_N), .QN(N404) );
  DFFRX1TF \id_ir_reg[3]  ( .D(N524), .CK(CLK), .RN(RST_N), .QN(N400) );
  DFFRX1TF \id_ir_reg[6]  ( .D(N521), .CK(CLK), .RN(RST_N), .QN(N403) );
  DFFRX1TF \id_ir_reg[5]  ( .D(N522), .CK(CLK), .RN(RST_N), .QN(N402) );
  DFFRX1TF \gr_reg[0][15]  ( .D(N953), .CK(CLK), .RN(RST_N), .QN(N677) );
  DFFRX1TF \gr_reg[0][14]  ( .D(N954), .CK(CLK), .RN(RST_N), .QN(N678) );
  DFFRX1TF \gr_reg[0][13]  ( .D(N955), .CK(CLK), .RN(RST_N), .QN(N679) );
  DFFRX1TF \gr_reg[4][15]  ( .D(N1001), .CK(CLK), .RN(RST_N), .QN(N613) );
  DFFRX1TF \gr_reg[4][14]  ( .D(N922), .CK(CLK), .RN(RST_N), .QN(N614) );
  DFFRX1TF \gr_reg[4][13]  ( .D(N923), .CK(CLK), .RN(RST_N), .QN(N615) );
  DFFRX1TF \gr_reg[2][15]  ( .D(N937), .CK(CLK), .RN(RST_N), .QN(N645) );
  DFFRX1TF \gr_reg[2][14]  ( .D(N938), .CK(CLK), .RN(RST_N), .QN(N646) );
  DFFRX1TF \gr_reg[2][13]  ( .D(N939), .CK(CLK), .RN(RST_N), .QN(N647) );
  DFFRX1TF \gr_reg[1][15]  ( .D(N945), .CK(CLK), .RN(RST_N), .QN(N661) );
  DFFRX1TF \gr_reg[1][14]  ( .D(N946), .CK(CLK), .RN(RST_N), .QN(N662) );
  DFFRX1TF \gr_reg[1][13]  ( .D(N947), .CK(CLK), .RN(RST_N), .QN(N663) );
  DFFRX1TF \gr_reg[0][12]  ( .D(N956), .CK(CLK), .RN(RST_N), .QN(N680) );
  DFFRX1TF \gr_reg[0][11]  ( .D(N957), .CK(CLK), .RN(RST_N), .QN(N681) );
  DFFRX1TF \gr_reg[0][10]  ( .D(N958), .CK(CLK), .RN(RST_N), .QN(N682) );
  DFFRX1TF \gr_reg[0][9]  ( .D(N959), .CK(CLK), .RN(RST_N), .QN(N683) );
  DFFRX1TF \gr_reg[0][8]  ( .D(N960), .CK(CLK), .RN(RST_N), .QN(N684) );
  DFFRX1TF \gr_reg[0][4]  ( .D(N996), .CK(CLK), .RN(RST_N), .QN(N688) );
  DFFRX1TF \gr_reg[0][3]  ( .D(N997), .CK(CLK), .RN(RST_N), .QN(N689) );
  DFFRX1TF \gr_reg[0][2]  ( .D(N998), .CK(CLK), .RN(RST_N), .QN(N690) );
  DFFRX1TF \gr_reg[0][1]  ( .D(N999), .CK(CLK), .RN(RST_N), .QN(N691) );
  DFFRX1TF \gr_reg[0][0]  ( .D(N1000), .CK(CLK), .RN(RST_N), .QN(N692) );
  DFFRX1TF \gr_reg[4][12]  ( .D(N924), .CK(CLK), .RN(RST_N), .QN(N6160) );
  DFFRX1TF \gr_reg[4][11]  ( .D(N925), .CK(CLK), .RN(RST_N), .QN(N617) );
  DFFRX1TF \gr_reg[4][10]  ( .D(N926), .CK(CLK), .RN(RST_N), .QN(N618) );
  DFFRX1TF \gr_reg[0][7]  ( .D(N993), .CK(CLK), .RN(RST_N), .QN(N685) );
  DFFRX1TF \gr_reg[0][6]  ( .D(N994), .CK(CLK), .RN(RST_N), .QN(N686) );
  DFFRX1TF \gr_reg[0][5]  ( .D(N995), .CK(CLK), .RN(RST_N), .QN(N687) );
  DFFRX1TF \gr_reg[1][12]  ( .D(N948), .CK(CLK), .RN(RST_N), .QN(N664) );
  DFFRX1TF \gr_reg[1][11]  ( .D(N949), .CK(CLK), .RN(RST_N), .QN(N665) );
  DFFRX1TF \gr_reg[1][10]  ( .D(N950), .CK(CLK), .RN(RST_N), .QN(N666) );
  DFFRX1TF \gr_reg[1][9]  ( .D(N951), .CK(CLK), .RN(RST_N), .QN(N667) );
  DFFRX1TF \gr_reg[1][8]  ( .D(N952), .CK(CLK), .RN(RST_N), .QN(N668) );
  DFFRX1TF \gr_reg[1][7]  ( .D(N985), .CK(CLK), .RN(RST_N), .QN(N669) );
  DFFRX1TF cf_reg ( .D(N5180), .CK(CLK), .RN(RST_N), .Q(CF) );
  DFFRX1TF \reg_A_reg[3]  ( .D(N4790), .CK(CLK), .RN(RST_N), .Q(REG_A[3]), 
        .QN(N1092) );
  DFFRX1TF \reg_A_reg[5]  ( .D(N444), .CK(CLK), .RN(RST_N), .Q(REG_A[5]), .QN(
        N836) );
  DFFRX2TF \id_ir_reg[9]  ( .D(N534), .CK(CLK), .RN(RST_N), .Q(N724), .QN(N571) );
  DFFRX2TF \reg_A_reg[14]  ( .D(N4830), .CK(CLK), .RN(RST_N), .Q(REG_A[14]), 
        .QN(N1101) );
  DFFNSRX2TF \reg_C_reg[2]  ( .D(N464), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[3]) );
  DFFNSRX2TF \reg_C_reg[4]  ( .D(N455), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[5]) );
  DFFNSRX2TF \reg_C_reg[6]  ( .D(N451), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[7]) );
  DFFNSRX2TF \reg_C_reg[5]  ( .D(N447), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[6]) );
  DFFNSRX2TF \reg_C_reg[3]  ( .D(N4820), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[4]) );
  DFFNSRX2TF \reg_C_reg[1]  ( .D(N491), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[2]) );
  DFFNSRX2TF \reg_C_reg[0]  ( .D(N500), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[1]) );
  DFFNSRX2TF \reg_C_reg[7]  ( .D(N5130), .CKN(CLK), .SN(1'b1), .RN(1'b1), .Q(
        D_ADDR[8]) );
  DFFRX2TF \reg_B_reg[0]  ( .D(N496), .CK(CLK), .RN(RST_N), .Q(REG_B[0]), .QN(
        N1130) );
  DFFRX2TF \reg_B_reg[2]  ( .D(N460), .CK(CLK), .RN(RST_N), .Q(REG_B[2]), .QN(
        N201) );
  DFFRX2TF \id_ir_reg[12]  ( .D(N531), .CK(CLK), .RN(RST_N), .Q(N223), .QN(N24) );
  ADDFHX2TF U3 ( .A(REG_A[1]), .B(REG_B[1]), .CI(ADD_X_285_3_N16), .CO(
        ADD_X_285_3_N15), .S(N471) );
  OAI21X4TF U4 ( .A0(N370), .A1(N126), .B0(N369), .Y(N500) );
  XOR2X4TF U5 ( .A(N365), .B(N364), .Y(N370) );
  ADDFHX4TF U6 ( .A(N406), .B(REG_A[6]), .CI(SUB_X_285_4_N11), .CO(
        SUB_X_285_4_N10), .S(N510) );
  ADDFX2TF U7 ( .A(N424), .B(REG_A[5]), .CI(SUB_X_285_4_N12), .CO(
        SUB_X_285_4_N11), .S(N509) );
  ADDFHX4TF U8 ( .A(N200), .B(REG_A[1]), .CI(SUB_X_285_4_N16), .CO(
        SUB_X_285_4_N15), .S(N505) );
  OAI222X2TF U9 ( .A0(N127), .A1(N362), .B0(N126), .B1(N384), .C0(N414), .C1(
        N217), .Y(N495) );
  AOI211X4TF U10 ( .A0(N519), .A1(N218), .B0(N6), .C0(N270), .Y(N7) );
  NAND2X1TF U11 ( .A(N387), .B(N204), .Y(N316) );
  INVX2TF U12 ( .A(N389), .Y(N121) );
  OAI211X1TF U13 ( .A0(N124), .A1(N194), .B0(N758), .C0(N762), .Y(N1) );
  OR2X1TF U14 ( .A(N742), .B(N1), .Y(N752) );
  NOR4BX1TF U15 ( .AN(N454), .B(N446), .C(N450), .D(N258), .Y(N2) );
  OAI2BB1X1TF U16 ( .A0N(N518), .A1N(N863), .B0(N2), .Y(N3) );
  AOI21X2TF U17 ( .A0(N337), .A1(N484), .B0(N3), .Y(N384) );
  AOI2BB2X1TF U18 ( .B0(N1174), .B1(IO_DATAINA[10]), .A0N(N361), .A1N(N125), 
        .Y(N4) );
  AOI22X1TF U19 ( .A0(N1172), .A1(REG_C[10]), .B0(N378), .B1(IO_DATAINB[10]), 
        .Y(N5) );
  OAI211X1TF U20 ( .A0(N371), .A1(N128), .B0(N4), .C0(N5), .Y(N4770) );
  AOI21X1TF U21 ( .A0(N134), .A1(N260), .B0(N412), .Y(N6) );
  OAI2BB1X4TF U22 ( .A0N(N337), .A1N(N485), .B0(N7), .Y(N365) );
  AOI2BB2X1TF U23 ( .B0(N1174), .B1(IO_DATAINA[11]), .A0N(N371), .A1N(N125), 
        .Y(N8) );
  AOI22X1TF U24 ( .A0(N1172), .A1(REG_C[11]), .B0(N220), .B1(IO_DATAINB[11]), 
        .Y(N9) );
  OAI211X1TF U25 ( .A0(N372), .A1(N128), .B0(N8), .C0(N9), .Y(N5100) );
  OAI21X1TF U26 ( .A0(N124), .A1(N202), .B0(N824), .Y(N10) );
  NOR3X1TF U27 ( .A(N822), .B(N823), .C(N10), .Y(N843) );
  AOI2BB2X1TF U28 ( .B0(N1174), .B1(IO_DATAINA[12]), .A0N(N372), .A1N(N125), 
        .Y(N11) );
  AOI22X1TF U29 ( .A0(N1172), .A1(REG_C[12]), .B0(N220), .B1(IO_DATAINB[12]), 
        .Y(N12) );
  OAI211XLTF U30 ( .A0(N385), .A1(N128), .B0(N11), .C0(N12), .Y(N5050) );
  AOI2BB1X1TF U31 ( .A0N(N124), .A1N(N831), .B0(N458), .Y(N295) );
  OAI21X1TF U32 ( .A0(N768), .A1(N176), .B0(N733), .Y(N13) );
  NOR3X1TF U33 ( .A(N731), .B(N732), .C(N13), .Y(N773) );
  AOI2BB2X1TF U34 ( .B0(N199), .B1(N1019), .A0N(N1023), .A1N(N1018), .Y(N140)
         );
  OA21XLTF U35 ( .A0(N696), .A1(I_ADDR[4]), .B0(N697), .Y(N14) );
  AOI222XLTF U36 ( .A0(I_ADDR[4]), .A1(N702), .B0(N709), .B1(D_ADDR[4]), .C0(
        N700), .C1(N14), .Y(N810) );
  CLKINVX1TF U37 ( .A(N218), .Y(N15) );
  OAI22X1TF U38 ( .A0(SUB_X_285_4_N1), .A1(N15), .B0(N16), .B1(N490), .Y(N589)
         );
  CLKINVX1TF U39 ( .A(N486), .Y(N16) );
  NAND2BX1TF U40 ( .AN(N876), .B(N921), .Y(N17) );
  OAI211X1TF U41 ( .A0(N1004), .A1(N392), .B0(N1003), .C0(N17), .Y(N1014) );
  OA21XLTF U42 ( .A0(N701), .A1(I_ADDR[6]), .B0(N706), .Y(N18) );
  AOI222XLTF U43 ( .A0(I_ADDR[6]), .A1(N702), .B0(N709), .B1(D_ADDR[6]), .C0(
        N700), .C1(N18), .Y(N808) );
  NOR4XLTF U44 ( .A(N1187), .B(N344), .C(N345), .D(N350), .Y(N19) );
  NAND4X1TF U45 ( .A(N19), .B(N374), .C(N379), .D(N381), .Y(N20) );
  NOR4XLTF U46 ( .A(N357), .B(N376), .C(N352), .D(N20), .Y(N21) );
  AND4X1TF U47 ( .A(N21), .B(N361), .C(N371), .D(N372), .Y(N22) );
  NAND4X1TF U48 ( .A(N22), .B(N385), .C(N386), .D(N384), .Y(N23) );
  OAI2BB2XLTF U49 ( .B0(N365), .B1(N23), .A0N(N1187), .A1N(ZF), .Y(N434) );
  OR2X2TF U50 ( .A(N1015), .B(N4850), .Y(N25) );
  OR3X1TF U51 ( .A(N1004), .B(N877), .C(N135), .Y(N867) );
  NOR2X4TF U52 ( .A(N200), .B(REG_B[0]), .Y(N26) );
  NOR2X1TF U53 ( .A(N200), .B(REG_B[0]), .Y(N787) );
  ADDFHX2TF U54 ( .A(REG_A[3]), .B(REG_B[3]), .CI(ADD_X_285_3_N14), .CO(
        ADD_X_285_3_N13), .S(N473) );
  CLKBUFX2TF U55 ( .A(N1180), .Y(N35) );
  INVX2TF U75 ( .A(N843), .Y(N849) );
  OR3X1TF U76 ( .A(N729), .B(N875), .C(N873), .Y(N1160) );
  INVX1TF U77 ( .A(N542), .Y(N237) );
  INVX2TF U78 ( .A(N223), .Y(N135) );
  XOR2X2TF U79 ( .A(N386), .B(N363), .Y(N364) );
  CLKXOR2X2TF U80 ( .A(N385), .B(N371), .Y(N363) );
  AO22X1TF U81 ( .A0(N1021), .A1(N1020), .B0(N401), .B1(N1019), .Y(N1167) );
  OAI22X1TF U82 ( .A0(N197), .A1(N1023), .B0(N1022), .B1(N403), .Y(N1166) );
  NAND4X2TF U83 ( .A(N198), .B(N185), .C(N180), .D(N885), .Y(N1176) );
  AND2X2TF U84 ( .A(N388), .B(N228), .Y(N1173) );
  OAI211XLTF U85 ( .A0(N1032), .A1(N1004), .B0(N540), .C0(N539), .Y(N541) );
  NAND2XLTF U86 ( .A(N392), .B(CODE_TYPE[3]), .Y(N878) );
  INVX2TF U87 ( .A(N723), .Y(N718) );
  ADDFX2TF U88 ( .A(N412), .B(REG_A[15]), .CI(SUB_X_285_4_N2), .CO(
        SUB_X_285_4_N1), .S(N519) );
  OA22X1TF U89 ( .A0(N381), .A1(N126), .B0(N382), .B1(N128), .Y(N1120) );
  AOI22X1TF U90 ( .A0(N579), .A1(N587), .B0(N667), .B1(N578), .Y(N951) );
  AOI22X1TF U91 ( .A0(N550), .A1(N564), .B0(N670), .B1(N549), .Y(N986) );
  AOI22X1TF U92 ( .A0(N552), .A1(N560), .B0(N658), .B1(N551), .Y(N982) );
  AOI22X1TF U93 ( .A0(N579), .A1(N5890), .B0(N665), .B1(N578), .Y(N949) );
  AOI22X1TF U94 ( .A0(N556), .A1(N566), .B0(N637), .B1(N555), .Y(N969) );
  AOI22X1TF U95 ( .A0(N585), .A1(N586), .B0(N636), .B1(N583), .Y(N936) );
  AOI22X1TF U96 ( .A0(N550), .A1(N566), .B0(N669), .B1(N549), .Y(N985) );
  AOI22X1TF U97 ( .A0(N556), .A1(N560), .B0(N642), .B1(N555), .Y(N974) );
  AOI22X1TF U98 ( .A0(N579), .A1(N586), .B0(N668), .B1(N578), .Y(N952) );
  AOI22X1TF U99 ( .A0(N552), .A1(N559), .B0(N659), .B1(N551), .Y(N983) );
  AOI22X1TF U100 ( .A0(N585), .A1(N587), .B0(N635), .B1(N583), .Y(N935) );
  AOI22X1TF U101 ( .A0(N581), .A1(N587), .B0(N651), .B1(N580), .Y(N943) );
  AOI22X1TF U102 ( .A0(N556), .A1(N564), .B0(N638), .B1(N555), .Y(N970) );
  AOI22X1TF U103 ( .A0(N581), .A1(N5880), .B0(N650), .B1(N580), .Y(N942) );
  AOI22X1TF U104 ( .A0(N585), .A1(N5890), .B0(N633), .B1(N583), .Y(N933) );
  AOI22X1TF U105 ( .A0(N581), .A1(N586), .B0(N652), .B1(N580), .Y(N944) );
  AOI22X1TF U106 ( .A0(N581), .A1(N5890), .B0(N649), .B1(N580), .Y(N941) );
  AOI22X1TF U107 ( .A0(N550), .A1(N559), .B0(N675), .B1(N549), .Y(N991) );
  AOI22X1TF U108 ( .A0(N585), .A1(N5880), .B0(N634), .B1(N583), .Y(N934) );
  AOI22X1TF U109 ( .A0(N556), .A1(N559), .B0(N643), .B1(N555), .Y(N975) );
  NOR4XLTF U110 ( .A(N817), .B(N333), .C(N818), .D(N332), .Y(N334) );
  AO22X1TF U111 ( .A0(N199), .A1(N1017), .B0(N1016), .B1(N1020), .Y(N1165) );
  OAI22X1TF U112 ( .A0(N678), .A1(N1660), .B0(N646), .B1(N163), .Y(N1105) );
  OAI22X1TF U113 ( .A0(N143), .A1(N600), .B0(N666), .B1(N160), .Y(N1086) );
  OAI22X1TF U114 ( .A0(N629), .A1(N1179), .B0(N661), .B1(N1178), .Y(N889) );
  OAI22X1TF U115 ( .A0(N682), .A1(N1660), .B0(N650), .B1(N163), .Y(N1085) );
  OAI22X1TF U116 ( .A0(N677), .A1(N1660), .B0(N645), .B1(N163), .Y(N1126) );
  OAI22X1TF U117 ( .A0(N144), .A1(N595), .B0(N661), .B1(N160), .Y(N1127) );
  OAI22X1TF U118 ( .A0(N631), .A1(N1179), .B0(N663), .B1(N1178), .Y(N901) );
  OAI22X1TF U119 ( .A0(N683), .A1(N1670), .B0(N651), .B1(N164), .Y(N1075) );
  OAI22X1TF U120 ( .A0(N680), .A1(N1670), .B0(N648), .B1(N164), .Y(N1149) );
  OAI22X1TF U121 ( .A0(N681), .A1(N1670), .B0(N649), .B1(N164), .Y(N1161) );
  OAI22X1TF U122 ( .A0(N679), .A1(N1670), .B0(N647), .B1(N164), .Y(N1069) );
  OAI22X1TF U123 ( .A0(N685), .A1(N1670), .B0(N653), .B1(N164), .Y(N725) );
  OAI22X1TF U124 ( .A0(N145), .A1(N602), .B0(N668), .B1(N160), .Y(N1052) );
  OAI22X1TF U125 ( .A0(N684), .A1(N1660), .B0(N652), .B1(N163), .Y(N1051) );
  OAI22X1TF U126 ( .A0(N687), .A1(N1670), .B0(N655), .B1(N164), .Y(N1027) );
  OAI22X1TF U127 ( .A0(N686), .A1(N1670), .B0(N654), .B1(N164), .Y(N1038) );
  OAI22X1TF U128 ( .A0(N688), .A1(N1660), .B0(N656), .B1(N163), .Y(N1044) );
  OAI22X1TF U129 ( .A0(N145), .A1(N606), .B0(N672), .B1(N160), .Y(N1045) );
  OAI22X1TF U130 ( .A0(N690), .A1(N1670), .B0(N658), .B1(N164), .Y(N1061) );
  OAI22X1TF U131 ( .A0(N691), .A1(N1660), .B0(N659), .B1(N163), .Y(N1116) );
  OAI22X1TF U132 ( .A0(N145), .A1(N607), .B0(N673), .B1(N160), .Y(N1097) );
  OAI22X1TF U133 ( .A0(N144), .A1(N610), .B0(N676), .B1(N160), .Y(N1139) );
  OAI22X1TF U134 ( .A0(N689), .A1(N1660), .B0(N657), .B1(N163), .Y(N1096) );
  OAI22X1TF U135 ( .A0(N692), .A1(N1660), .B0(N660), .B1(N163), .Y(N1138) );
  AND2X2TF U136 ( .A(N1010), .B(N1020), .Y(N1011) );
  NAND3XLTF U137 ( .A(N494), .B(N842), .C(N490), .Y(N588) );
  AND2X2TF U138 ( .A(\OPER1_R1[2] ), .B(N144), .Y(N156) );
  AND2X2TF U139 ( .A(N1010), .B(N143), .Y(N165) );
  AND2X2TF U140 ( .A(N1021), .B(N143), .Y(N162) );
  OAI31XLTF U141 ( .A0(IO_STATUS[0]), .A1(IO_STATUS[1]), .A2(N720), .B0(N719), 
        .Y(NEXT_STATE[1]) );
  AND2X2TF U142 ( .A(N1016), .B(N143), .Y(N159) );
  CLKBUFX2TF U143 ( .A(N570), .Y(N146) );
  AND2X2TF U144 ( .A(OPER3_R3[2]), .B(N885), .Y(N1186) );
  AND2X2TF U145 ( .A(N388), .B(N251), .Y(N1175) );
  AOI32X1TF U146 ( .A0(N542), .A1(N543), .A2(N391), .B0(N541), .B1(N543), .Y(
        N570) );
  INVX1TF U147 ( .A(N835), .Y(N763) );
  CLKINVX1TF U148 ( .A(N316), .Y(N303) );
  NAND2XLTF U149 ( .A(N393), .B(REG_A[5]), .Y(N757) );
  NAND3BXLTF U150 ( .AN(N882), .B(N1003), .C(N1004), .Y(N259) );
  ADDFHX2TF U151 ( .A(N423), .B(REG_A[4]), .CI(SUB_X_285_4_N13), .CO(
        SUB_X_285_4_N12), .S(N508) );
  CLKINVX2TF U152 ( .A(N388), .Y(N150) );
  ADDFHX2TF U153 ( .A(N204), .B(REG_A[3]), .CI(SUB_X_285_4_N14), .CO(
        SUB_X_285_4_N13), .S(N507) );
  OAI32X1TF U154 ( .A0(STATE[1]), .A1(STATE[3]), .A2(N554), .B0(N721), .B1(
        N183), .Y(N110) );
  OR2X1TF U155 ( .A(REG_B[2]), .B(N764), .Y(N203) );
  AOI22X1TF U156 ( .A0(N735), .A1(REG_A[0]), .B0(N787), .B1(REG_A[1]), .Y(N463) );
  NAND2XLTF U157 ( .A(N26), .B(REG_A[12]), .Y(N425) );
  NAND2XLTF U158 ( .A(N26), .B(REG_A[3]), .Y(N766) );
  AND2X2TF U159 ( .A(N200), .B(N1130), .Y(N821) );
  INVX2TF U160 ( .A(N1188), .Y(N149) );
  NAND2XLTF U161 ( .A(STATE[0]), .B(N183), .Y(N710) );
  NAND4XLTF U162 ( .A(N554), .B(N671), .C(N670), .D(N669), .Y(N713) );
  NAND2XLTF U163 ( .A(STATE[1]), .B(N179), .Y(N4810) );
  INVX2TF U164 ( .A(N867), .Y(N122) );
  INVX2TF U165 ( .A(N821), .Y(N123) );
  INVX2TF U166 ( .A(N821), .Y(N124) );
  INVX2TF U167 ( .A(N1175), .Y(N125) );
  INVX2TF U168 ( .A(N1175), .Y(N126) );
  INVX2TF U169 ( .A(N1173), .Y(N127) );
  INVX2TF U170 ( .A(N1173), .Y(N128) );
  INVX2TF U171 ( .A(N1047), .Y(N129) );
  INVX2TF U172 ( .A(N1047), .Y(N130) );
  INVX2TF U173 ( .A(N1165), .Y(N131) );
  INVX2TF U174 ( .A(N1165), .Y(N132) );
  INVX2TF U175 ( .A(N25), .Y(N133) );
  INVX2TF U176 ( .A(N25), .Y(N134) );
  INVX2TF U177 ( .A(N1166), .Y(N136) );
  INVX2TF U178 ( .A(N1166), .Y(N137) );
  INVX2TF U179 ( .A(N1167), .Y(N138) );
  INVX2TF U180 ( .A(N1167), .Y(N139) );
  INVX2TF U181 ( .A(N140), .Y(N141) );
  INVX2TF U182 ( .A(N140), .Y(N142) );
  INVX2TF U183 ( .A(N1160), .Y(N143) );
  INVX2TF U184 ( .A(N1160), .Y(N144) );
  INVX2TF U185 ( .A(N1160), .Y(N145) );
  AOI22XLTF U186 ( .A0(N307), .A1(N846), .B0(N740), .B1(N844), .Y(N262) );
  NOR3X2TF U187 ( .A(N724), .B(N210), .C(\OPER1_R1[2] ), .Y(N1010) );
  AOI22X2TF U188 ( .A0(REG_C[10]), .A1(N568), .B0(N573), .B1(D_DATAIN[2]), .Y(
        N5880) );
  AOI22X2TF U189 ( .A0(REG_C[11]), .A1(N568), .B0(N573), .B1(D_DATAIN[3]), .Y(
        N5890) );
  AOI22X2TF U190 ( .A0(REG_C[8]), .A1(N568), .B0(N573), .B1(D_DATAIN[0]), .Y(
        N586) );
  AOI22X2TF U191 ( .A0(REG_C[9]), .A1(N568), .B0(N573), .B1(D_DATAIN[1]), .Y(
        N587) );
  AOI22X2TF U192 ( .A0(D_ADDR[3]), .A1(N546), .B0(N545), .B1(D_DATAIN[2]), .Y(
        N560) );
  AOI22X2TF U193 ( .A0(D_ADDR[2]), .A1(N546), .B0(N545), .B1(D_DATAIN[1]), .Y(
        N559) );
  AOI22X2TF U194 ( .A0(D_ADDR[7]), .A1(N546), .B0(N545), .B1(D_DATAIN[6]), .Y(
        N564) );
  AOI22X2TF U195 ( .A0(D_ADDR[8]), .A1(N546), .B0(N545), .B1(D_DATAIN[7]), .Y(
        N566) );
  NOR2X4TF U196 ( .A(N200), .B(N1130), .Y(N735) );
  AOI32X1TF U197 ( .A0(N195), .A1(N205), .A2(N716), .B0(STATE[0]), .B1(N4810), 
        .Y(N166) );
  NOR3X4TF U198 ( .A(N857), .B(REG_B[3]), .C(REG_B[2]), .Y(N852) );
  NOR2BX2TF U199 ( .AN(CODE_TYPE[4]), .B(CODE_TYPE[3]), .Y(N391) );
  OAI22X2TF U200 ( .A0(N5160), .A1(N544), .B0(N721), .B1(N716), .Y(N703) );
  NOR3X4TF U201 ( .A(N572), .B(N571), .C(N553), .Y(N556) );
  NOR3X4TF U202 ( .A(N572), .B(N571), .C(N582), .Y(N585) );
  NOR3X4TF U203 ( .A(N571), .B(N210), .C(N582), .Y(N581) );
  OAI211XLTF U204 ( .A0(N723), .A1(N711), .B0(N710), .C0(N1191), .Y(
        NEXT_STATE[0]) );
  NOR3X4TF U205 ( .A(N195), .B(N205), .C(N723), .Y(N545) );
  NAND2X2TF U206 ( .A(N554), .B(STATE[1]), .Y(N723) );
  OAI22XLTF U207 ( .A0(N656), .A1(N1181), .B0(N423), .B1(N1180), .Y(N909) );
  OAI22XLTF U208 ( .A0(N657), .A1(N1181), .B0(N204), .B1(N1180), .Y(N1088) );
  OAI22XLTF U209 ( .A0(N654), .A1(N1181), .B0(N406), .B1(N1180), .Y(N913) );
  OAI22XLTF U210 ( .A0(N655), .A1(N1181), .B0(N424), .B1(N1180), .Y(N917) );
  OAI22XLTF U211 ( .A0(N658), .A1(N1181), .B0(N201), .B1(N1180), .Y(N1054) );
  OAI22XLTF U212 ( .A0(N659), .A1(N1181), .B0(N200), .B1(N1180), .Y(N1108) );
  INVX2TF U213 ( .A(N1186), .Y(N147) );
  INVX2TF U214 ( .A(N1186), .Y(N148) );
  INVX2TF U215 ( .A(N1191), .Y(N151) );
  INVX2TF U216 ( .A(N842), .Y(N152) );
  NOR2X1TF U217 ( .A(N1004), .B(N1030), .Y(N390) );
  CLKBUFX2TF U218 ( .A(N1171), .Y(N153) );
  CLKBUFX2TF U219 ( .A(N1163), .Y(N154) );
  NOR2BX2TF U220 ( .AN(N143), .B(N1018), .Y(N1163) );
  CLKBUFX2TF U221 ( .A(N1176), .Y(N155) );
  OAI31X4TF U222 ( .A0(N1015), .A1(N1014), .A2(N1013), .B0(N1012), .Y(N1047)
         );
  NOR2X2TF U223 ( .A(REG_B[3]), .B(N201), .Y(N848) );
  INVX2TF U224 ( .A(N156), .Y(N157) );
  INVX2TF U225 ( .A(N156), .Y(N158) );
  INVX2TF U226 ( .A(N159), .Y(N160) );
  INVX2TF U227 ( .A(N159), .Y(N161) );
  INVX2TF U228 ( .A(N162), .Y(N163) );
  INVX2TF U229 ( .A(N162), .Y(N164) );
  OAI21X2TF U230 ( .A0(N881), .A1(N908), .B0(N1012), .Y(N1129) );
  OAI211X1TF U231 ( .A0(CODE_TYPE[3]), .A1(N874), .B0(N1012), .C0(N182), .Y(
        N883) );
  INVX2TF U232 ( .A(N165), .Y(N1660) );
  INVX2TF U233 ( .A(N165), .Y(N1670) );
  CLKBUFX2TF U234 ( .A(N1179), .Y(N1680) );
  OAI22XLTF U235 ( .A0(N636), .A1(N1179), .B0(N668), .B1(N1178), .Y(N905) );
  OAI22XLTF U236 ( .A0(N635), .A1(N1179), .B0(N667), .B1(N1178), .Y(N897) );
  OAI22XLTF U237 ( .A0(N630), .A1(N1179), .B0(N662), .B1(N1178), .Y(N893) );
  NOR3X4TF U238 ( .A(N571), .B(N210), .C(N553), .Y(N552) );
  CLKBUFX2TF U239 ( .A(N1174), .Y(N169) );
  NOR2X1TF U240 ( .A(N223), .B(N1119), .Y(N1174) );
  AOI2BB2X2TF U241 ( .B0(D_DATAIN[5]), .B1(N573), .A0N(N421), .A1N(N146), .Y(
        N591) );
  AOI2BB2X2TF U242 ( .B0(D_DATAIN[6]), .B1(N573), .A0N(N416), .A1N(N146), .Y(
        N593) );
  AOI2BB2X2TF U243 ( .B0(D_DATAIN[7]), .B1(N573), .A0N(N414), .A1N(N146), .Y(
        N584) );
  AOI22X2TF U244 ( .A0(REG_C[12]), .A1(N568), .B0(N573), .B1(D_DATAIN[4]), .Y(
        N590) );
  NOR3X4TF U245 ( .A(N186), .B(N875), .C(N876), .Y(N573) );
  AOI22X2TF U246 ( .A0(D_ADDR[1]), .A1(N546), .B0(N545), .B1(D_DATAIN[0]), .Y(
        N558) );
  AOI22X2TF U247 ( .A0(D_ADDR[6]), .A1(N546), .B0(N545), .B1(D_DATAIN[5]), .Y(
        N563) );
  AOI22X2TF U248 ( .A0(D_ADDR[5]), .A1(N546), .B0(N545), .B1(D_DATAIN[4]), .Y(
        N562) );
  AOI22X2TF U249 ( .A0(D_ADDR[4]), .A1(N546), .B0(N545), .B1(D_DATAIN[3]), .Y(
        N561) );
  NOR3X4TF U250 ( .A(N195), .B(N723), .C(STATE[0]), .Y(N546) );
  AOI22XLTF U251 ( .A0(N735), .A1(REG_A[13]), .B0(N787), .B1(REG_A[12]), .Y(
        N736) );
  CMPR32X2TF U252 ( .A(REG_A[15]), .B(REG_B[15]), .C(ADD_X_285_3_N2), .CO(N486), .S(N485) );
  CMPR22X2TF U253 ( .A(REG_B[0]), .B(REG_A[0]), .CO(ADD_X_285_3_N16), .S(N470)
         );
  XOR2X1TF U254 ( .A(REG_A[0]), .B(REG_B[0]), .Y(N504) );
  NAND2BX4TF U255 ( .AN(REG_A[0]), .B(REG_B[0]), .Y(SUB_X_285_4_N16) );
  CLKINVX6TF U256 ( .A(N365), .Y(N362) );
  NOR2X4TF U257 ( .A(N1004), .B(N880), .Y(N389) );
  NOR2X2TF U258 ( .A(N181), .B(N186), .Y(N1032) );
  AOI21X1TF U259 ( .A0(N480), .A1(N219), .B0(N282), .Y(N371) );
  INVX2TF U260 ( .A(N123), .Y(N393) );
  AO21X1TF U261 ( .A0(IO_DATAINA[9]), .A1(N169), .B0(N360), .Y(N4720) );
  AOI21X2TF U262 ( .A0(N482), .A1(N219), .B0(N257), .Y(N385) );
  CLKBUFX2TF U263 ( .A(N337), .Y(N219) );
  NAND2X1TF U264 ( .A(N181), .B(N223), .Y(N876) );
  OAI2BB1X1TF U265 ( .A0N(N219), .A1N(N478), .B0(N336), .Y(N357) );
  AOI21X2TF U266 ( .A0(N483), .A1(N337), .B0(N250), .Y(N386) );
  NOR3X1TF U267 ( .A(N569), .B(N223), .C(N181), .Y(N874) );
  AOI211XLTF U268 ( .A0(STATE[0]), .A1(N718), .B0(N217), .C0(N717), .Y(N719)
         );
  AOI31X1TF U269 ( .A0(N135), .A1(N392), .A2(N921), .B0(N544), .Y(N715) );
  NAND2X1TF U270 ( .A(N576), .B(N197), .Y(N582) );
  NAND2X1TF U271 ( .A(N197), .B(N557), .Y(N553) );
  OAI2BB2X1TF U272 ( .B0(N544), .B1(N146), .A0N(N573), .A1N(N545), .Y(N557) );
  CLKBUFX2TF U273 ( .A(N388), .Y(N217) );
  CLKBUFX2TF U274 ( .A(N863), .Y(N218) );
  NAND2X1TF U275 ( .A(N1012), .B(N1013), .Y(N1023) );
  NOR2X1TF U276 ( .A(N883), .B(N908), .Y(N885) );
  NAND3X2TF U277 ( .A(N883), .B(N1129), .C(N1152), .Y(N1180) );
  AOI21X1TF U278 ( .A0(N543), .A1(N146), .B0(N544), .Y(N576) );
  INVX2TF U279 ( .A(N388), .Y(N1172) );
  INVX2TF U280 ( .A(N861), .Y(N430) );
  NOR2X2TF U281 ( .A(CODE_TYPE[3]), .B(CODE_TYPE[4]), .Y(N921) );
  NAND2X1TF U282 ( .A(N181), .B(N186), .Y(N1009) );
  OR2X2TF U283 ( .A(N240), .B(N239), .Y(N337) );
  NOR2X2TF U284 ( .A(N135), .B(N569), .Y(N542) );
  OAI211XLTF U285 ( .A0(IO_CONTROL[4]), .A1(N713), .B0(N712), .C0(STATE[1]), 
        .Y(N720) );
  AOI22XLTF U286 ( .A0(REG_A[5]), .A1(N1047), .B0(IO_CONTROL[5]), .B1(N1165), 
        .Y(N1026) );
  NAND2X1TF U287 ( .A(N1012), .B(N1014), .Y(N1022) );
  NAND2X1TF U288 ( .A(N259), .B(N217), .Y(N1187) );
  NAND3X2TF U289 ( .A(OPER3_R3[0]), .B(OPER3_R3[1]), .C(N885), .Y(N1179) );
  INVX2TF U290 ( .A(N873), .Y(N1012) );
  INVX2TF U291 ( .A(N1191), .Y(N1193) );
  NAND3X1TF U292 ( .A(N179), .B(N183), .C(N712), .Y(N1191) );
  INVX2TF U293 ( .A(N1188), .Y(N1189) );
  NOR2X2TF U294 ( .A(N577), .B(N582), .Y(N579) );
  NOR2X2TF U295 ( .A(N577), .B(N553), .Y(N550) );
  NOR2X1TF U296 ( .A(N724), .B(N572), .Y(N1016) );
  INVX2TF U297 ( .A(N546), .Y(N544) );
  INVX2TF U298 ( .A(N921), .Y(N875) );
  NAND2X2TF U299 ( .A(N864), .B(N848), .Y(N828) );
  NAND3X1TF U300 ( .A(N391), .B(N1032), .C(N217), .Y(N1119) );
  NAND3X2TF U301 ( .A(N223), .B(N1032), .C(N921), .Y(N857) );
  NAND2X2TF U302 ( .A(CODE_TYPE[2]), .B(N542), .Y(N880) );
  NOR2X1TF U303 ( .A(N191), .B(N182), .Y(N1006) );
  AND2X2TF U304 ( .A(N554), .B(N226), .Y(N388) );
  NOR3BX1TF U305 ( .AN(STATE[0]), .B(STATE[3]), .C(STATE[1]), .Y(N226) );
  OAI32XLTF U306 ( .A0(N205), .A1(STATE[1]), .A2(N554), .B0(N723), .B1(N205), 
        .Y(NEXT_STATE[3]) );
  NOR2XLTF U307 ( .A(STATE[1]), .B(N179), .Y(N722) );
  AO22X1TF U308 ( .A0(N383), .A1(CF_BUF), .B0(N1187), .B1(CF), .Y(N5180) );
  AOI22XLTF U309 ( .A0(REG_A[6]), .A1(N1047), .B0(IO_CONTROL[6]), .B1(N1165), 
        .Y(N1037) );
  NOR2BX1TF U310 ( .AN(N402), .B(N1022), .Y(N1017) );
  NAND2X1TF U311 ( .A(N705), .B(I_ADDR[8]), .Y(N714) );
  NOR2X1TF U312 ( .A(N706), .B(N212), .Y(N705) );
  OAI2BB2XLTF U313 ( .B0(N1193), .B1(N135), .A0N(N1193), .A1N(I_DATAIN[4]), 
        .Y(N531) );
  OAI2BB2XLTF U314 ( .B0(N1189), .B1(N185), .A0N(N1189), .A1N(I_DATAIN[1]), 
        .Y(N526) );
  OAI2BB2XLTF U315 ( .B0(N1193), .B1(N181), .A0N(N1193), .A1N(I_DATAIN[5]), 
        .Y(N530) );
  OAI2BB2XLTF U316 ( .B0(N1189), .B1(N402), .A0N(N1189), .A1N(I_DATAIN[5]), 
        .Y(N522) );
  OAI2BB2XLTF U317 ( .B0(N1189), .B1(N180), .A0N(N1189), .A1N(I_DATAIN[2]), 
        .Y(N525) );
  OAI2BB2XLTF U318 ( .B0(N1193), .B1(N191), .A0N(N1193), .A1N(I_DATAIN[6]), 
        .Y(N529) );
  OAI2BB2XLTF U319 ( .B0(N1193), .B1(N571), .A0N(N1193), .A1N(I_DATAIN[1]), 
        .Y(N534) );
  OAI2BB2XLTF U320 ( .B0(N1189), .B1(N198), .A0N(N1189), .A1N(I_DATAIN[0]), 
        .Y(N527) );
  OAI2BB2XLTF U321 ( .B0(N1193), .B1(N572), .A0N(N151), .A1N(I_DATAIN[0]), .Y(
        N535) );
  OAI2BB2XLTF U322 ( .B0(N1193), .B1(N197), .A0N(N151), .A1N(I_DATAIN[2]), .Y(
        N533) );
  OAI2BB2XLTF U323 ( .B0(N1189), .B1(N403), .A0N(N149), .A1N(I_DATAIN[6]), .Y(
        N521) );
  NAND4X1TF U324 ( .A(N195), .B(N179), .C(N183), .D(STATE[0]), .Y(N1188) );
  INVX2TF U325 ( .A(N579), .Y(N578) );
  INVX2TF U326 ( .A(N585), .Y(N583) );
  INVX2TF U327 ( .A(N581), .Y(N580) );
  INVX2TF U328 ( .A(N556), .Y(N555) );
  INVX2TF U329 ( .A(N592), .Y(N594) );
  NAND2X2TF U330 ( .A(N557), .B(N1010), .Y(N547) );
  INVX2TF U331 ( .A(N552), .Y(N551) );
  INVX2TF U332 ( .A(N565), .Y(N567) );
  OAI221XLTF U333 ( .A0(N718), .A1(N538), .B0(N723), .B1(N721), .C0(N537), .Y(
        N1002) );
  NAND4X1TF U334 ( .A(N179), .B(N183), .C(STATE[0]), .D(STATE[3]), .Y(N873) );
  NOR2X1TF U335 ( .A(STATE[3]), .B(STATE[0]), .Y(N712) );
  OAI221XLTF U336 ( .A0(REG_A[2]), .A1(N121), .B0(N177), .B1(N842), .C0(N134), 
        .Y(N781) );
  OAI221XLTF U337 ( .A0(REG_A[1]), .A1(N121), .B0(N1112), .B1(N842), .C0(N134), 
        .Y(N772) );
  INVX2TF U338 ( .A(N390), .Y(N842) );
  NAND2X1TF U339 ( .A(N26), .B(REG_A[10]), .Y(N806) );
  NAND2X1TF U340 ( .A(N26), .B(REG_A[11]), .Y(N760) );
  NAND2X1TF U341 ( .A(N26), .B(REG_A[7]), .Y(N756) );
  NAND2X1TF U342 ( .A(N26), .B(REG_A[8]), .Y(N733) );
  NAND2X1TF U343 ( .A(N921), .B(N874), .Y(N396) );
  NAND2BX1TF U344 ( .AN(N1004), .B(N230), .Y(N490) );
  NAND2X1TF U345 ( .A(N181), .B(N135), .Y(N1005) );
  NOR3X1TF U346 ( .A(N225), .B(N4850), .C(N863), .Y(N494) );
  OAI21X1TF U347 ( .A0(N722), .A1(N721), .B0(N1188), .Y(NEXT_STATE[2]) );
  INVX2TF U348 ( .A(N1187), .Y(N383) );
  OAI21X1TF U349 ( .A0(N624), .A1(N157), .B0(N1046), .Y(N453) );
  AOI211X1TF U350 ( .A0(N1163), .A1(IO_DATAOUTB[4]), .B0(N1045), .C0(N1044), 
        .Y(N1046) );
  OAI21X1TF U351 ( .A0(N625), .A1(N157), .B0(N1098), .Y(N4800) );
  AOI211X1TF U352 ( .A0(N1163), .A1(IO_DATAOUTB[3]), .B0(N1097), .C0(N1096), 
        .Y(N1098) );
  OAI21X1TF U353 ( .A0(N613), .A1(N157), .B0(N1128), .Y(N493) );
  AOI211X1TF U354 ( .A0(N1163), .A1(N216), .B0(N1127), .C0(N1126), .Y(N1128)
         );
  OAI21X1TF U355 ( .A0(N620), .A1(N157), .B0(N1053), .Y(N457) );
  AOI211X1TF U356 ( .A0(N1163), .A1(IO_DATAOUTB[8]), .B0(N1052), .C0(N1051), 
        .Y(N1053) );
  OAI21X1TF U357 ( .A0(N628), .A1(N157), .B0(N1140), .Y(N498) );
  AOI211X1TF U358 ( .A0(N1163), .A1(IO_DATAOUTB[0]), .B0(N1139), .C0(N1138), 
        .Y(N1140) );
  OAI21X1TF U359 ( .A0(N618), .A1(N157), .B0(N1087), .Y(N4750) );
  AOI211X1TF U360 ( .A0(N1163), .A1(IO_DATAOUTB[10]), .B0(N1086), .C0(N1085), 
        .Y(N1087) );
  OAI21X1TF U361 ( .A0(N627), .A1(N157), .B0(N1118), .Y(N489) );
  AOI211X1TF U362 ( .A0(N1163), .A1(IO_DATAOUTB[1]), .B0(N1117), .C0(N1116), 
        .Y(N1118) );
  OAI22X1TF U363 ( .A0(N145), .A1(N609), .B0(N675), .B1(N161), .Y(N1117) );
  OAI21X1TF U364 ( .A0(N614), .A1(N157), .B0(N1107), .Y(N4840) );
  AOI211X1TF U365 ( .A0(N154), .A1(N215), .B0(N1106), .C0(N1105), .Y(N1107) );
  OAI22X1TF U366 ( .A0(N144), .A1(N596), .B0(N662), .B1(N161), .Y(N1106) );
  OAI21X1TF U367 ( .A0(N622), .A1(N158), .B0(N1040), .Y(N449) );
  AOI211X1TF U368 ( .A0(N154), .A1(IO_DATAOUTB[6]), .B0(N1039), .C0(N1038), 
        .Y(N1040) );
  OAI22X1TF U369 ( .A0(N145), .A1(N604), .B0(N670), .B1(N161), .Y(N1039) );
  OAI21X1TF U370 ( .A0(N621), .A1(N158), .B0(N727), .Y(N433) );
  AOI211X1TF U371 ( .A0(N154), .A1(IO_DATAOUTB[7]), .B0(N726), .C0(N725), .Y(
        N727) );
  OAI22X1TF U372 ( .A0(N144), .A1(N603), .B0(N669), .B1(N161), .Y(N726) );
  OAI21X1TF U373 ( .A0(N615), .A1(N158), .B0(N1071), .Y(N466) );
  AOI211X1TF U374 ( .A0(N154), .A1(N214), .B0(N1070), .C0(N1069), .Y(N1071) );
  OAI22X1TF U375 ( .A0(N145), .A1(N597), .B0(N663), .B1(N161), .Y(N1070) );
  OAI21X1TF U376 ( .A0(N619), .A1(N158), .B0(N1077), .Y(N4700) );
  AOI211X1TF U377 ( .A0(N154), .A1(IO_DATAOUTB[9]), .B0(N1076), .C0(N1075), 
        .Y(N1077) );
  OAI22X1TF U378 ( .A0(N144), .A1(N601), .B0(N667), .B1(N161), .Y(N1076) );
  OAI21X1TF U379 ( .A0(N623), .A1(N158), .B0(N1029), .Y(N445) );
  AOI211X1TF U380 ( .A0(N154), .A1(IO_DATAOUTB[5]), .B0(N1028), .C0(N1027), 
        .Y(N1029) );
  OAI22X1TF U381 ( .A0(N145), .A1(N605), .B0(N671), .B1(N161), .Y(N1028) );
  OAI21X1TF U382 ( .A0(N6160), .A1(N158), .B0(N1151), .Y(N503) );
  AOI211X1TF U383 ( .A0(N154), .A1(IO_DATAOUTB[12]), .B0(N1150), .C0(N1149), 
        .Y(N1151) );
  OAI22X1TF U384 ( .A0(N144), .A1(N598), .B0(N664), .B1(N161), .Y(N1150) );
  OAI21X1TF U385 ( .A0(N617), .A1(N158), .B0(N1164), .Y(N5080) );
  AOI211X1TF U386 ( .A0(N154), .A1(IO_DATAOUTB[11]), .B0(N1162), .C0(N1161), 
        .Y(N1164) );
  OAI22X1TF U387 ( .A0(N145), .A1(N599), .B0(N665), .B1(N161), .Y(N1162) );
  OAI21X1TF U388 ( .A0(N626), .A1(N158), .B0(N1063), .Y(N462) );
  AOI211X1TF U389 ( .A0(N154), .A1(IO_DATAOUTB[2]), .B0(N1062), .C0(N1061), 
        .Y(N1063) );
  OAI22X1TF U390 ( .A0(N144), .A1(N608), .B0(N674), .B1(N161), .Y(N1062) );
  OAI21X1TF U391 ( .A0(N1171), .A1(N680), .B0(N1148), .Y(N502) );
  AOI211X1TF U392 ( .A0(IO_DATAOUTB[12]), .A1(N141), .B0(N1147), .C0(N1146), 
        .Y(N1148) );
  OAI21X1TF U393 ( .A0(N1171), .A1(N681), .B0(N1159), .Y(N5070) );
  AOI211X1TF U394 ( .A0(IO_DATAOUTB[11]), .A1(N141), .B0(N1158), .C0(N1157), 
        .Y(N1159) );
  OAI21X1TF U395 ( .A0(N1171), .A1(N677), .B0(N1125), .Y(N492) );
  AOI211X1TF U396 ( .A0(N216), .A1(N141), .B0(N1124), .C0(N1123), .Y(N1125) );
  OAI21X1TF U397 ( .A0(N1171), .A1(N684), .B0(N1050), .Y(N456) );
  AOI211X1TF U398 ( .A0(IO_DATAOUTB[8]), .A1(N141), .B0(N1049), .C0(N1048), 
        .Y(N1050) );
  OAI21X1TF U399 ( .A0(N153), .A1(N690), .B0(N1060), .Y(N461) );
  AOI211X1TF U400 ( .A0(IO_DATAOUTB[2]), .A1(N142), .B0(N1059), .C0(N1058), 
        .Y(N1060) );
  OAI21X1TF U401 ( .A0(N1171), .A1(N682), .B0(N1084), .Y(N4740) );
  AOI211X1TF U402 ( .A0(IO_DATAOUTB[10]), .A1(N142), .B0(N1083), .C0(N1082), 
        .Y(N1084) );
  OAI21X1TF U403 ( .A0(N1171), .A1(N683), .B0(N1074), .Y(N469) );
  AOI211X1TF U404 ( .A0(IO_DATAOUTB[9]), .A1(N142), .B0(N1073), .C0(N1072), 
        .Y(N1074) );
  OAI21X1TF U405 ( .A0(N153), .A1(N685), .B0(N1170), .Y(N5110) );
  AOI211X1TF U406 ( .A0(IO_DATAOUTB[7]), .A1(N141), .B0(N1169), .C0(N1168), 
        .Y(N1170) );
  OAI21X1TF U407 ( .A0(N153), .A1(N679), .B0(N1068), .Y(N465) );
  AOI211X1TF U408 ( .A0(N214), .A1(N141), .B0(N1067), .C0(N1066), .Y(N1068) );
  OAI21X1TF U409 ( .A0(N153), .A1(N678), .B0(N1104), .Y(N4830) );
  AOI211X1TF U410 ( .A0(N215), .A1(N141), .B0(N1103), .C0(N1102), .Y(N1104) );
  OAI21X1TF U411 ( .A0(N153), .A1(N689), .B0(N1095), .Y(N4790) );
  AOI211X1TF U412 ( .A0(IO_DATAOUTB[3]), .A1(N141), .B0(N1094), .C0(N1093), 
        .Y(N1095) );
  OAI21X1TF U413 ( .A0(N153), .A1(N691), .B0(N1115), .Y(N488) );
  AOI211X1TF U414 ( .A0(IO_DATAOUTB[1]), .A1(N142), .B0(N1114), .C0(N1113), 
        .Y(N1115) );
  OAI21X1TF U415 ( .A0(N153), .A1(N692), .B0(N1137), .Y(N497) );
  AOI211X1TF U416 ( .A0(IO_DATAOUTB[0]), .A1(N142), .B0(N1136), .C0(N1135), 
        .Y(N1137) );
  OAI21X1TF U417 ( .A0(N624), .A1(N148), .B0(N912), .Y(N441) );
  NOR3X1TF U418 ( .A(N911), .B(N910), .C(N909), .Y(N912) );
  OAI22X1TF U419 ( .A0(N640), .A1(N1680), .B0(N672), .B1(N1178), .Y(N910) );
  OAI22X1TF U420 ( .A0(N688), .A1(N155), .B0(N401), .B1(N1177), .Y(N911) );
  OAI211X1TF U421 ( .A0(N1171), .A1(N687), .B0(N1026), .C0(N1025), .Y(N444) );
  AOI21X1TF U422 ( .A0(IO_DATAOUTB[5]), .A1(N142), .B0(N1024), .Y(N1025) );
  OAI211X1TF U423 ( .A0(N1171), .A1(N686), .B0(N1037), .C0(N1036), .Y(N448) );
  AOI21X1TF U424 ( .A0(IO_DATAOUTB[6]), .A1(N142), .B0(N1035), .Y(N1036) );
  OAI211X1TF U425 ( .A0(N1171), .A1(N688), .B0(N1043), .C0(N1042), .Y(N452) );
  AOI21X1TF U426 ( .A0(IO_DATAOUTB[4]), .A1(N142), .B0(N1041), .Y(N1042) );
  NOR2X1TF U427 ( .A(N571), .B(N210), .Y(N1021) );
  NOR2X1TF U428 ( .A(N1022), .B(N402), .Y(N1019) );
  AOI22X1TF U429 ( .A0(REG_A[4]), .A1(N1047), .B0(IO_CONTROL[4]), .B1(N1165), 
        .Y(N1043) );
  AOI31X4TF U430 ( .A0(N403), .A1(N401), .A2(N1017), .B0(N1011), .Y(N1171) );
  INVX2TF U431 ( .A(N1023), .Y(N1020) );
  OAI211X1TF U432 ( .A0(N191), .A1(N1009), .B0(N1008), .C0(N1007), .Y(N1013)
         );
  AOI32X1TF U433 ( .A0(N391), .A1(N230), .A2(N569), .B0(N1006), .B1(N1005), 
        .Y(N1008) );
  OAI21X1TF U434 ( .A0(N627), .A1(N148), .B0(N1111), .Y(N487) );
  NOR3X1TF U435 ( .A(N1110), .B(N1109), .C(N1108), .Y(N1111) );
  OAI22X1TF U436 ( .A0(N643), .A1(N1179), .B0(N675), .B1(N221), .Y(N1109) );
  OAI22X1TF U437 ( .A0(N691), .A1(N1176), .B0(N185), .B1(N1129), .Y(N1110) );
  OAI21X1TF U438 ( .A0(N626), .A1(N148), .B0(N1057), .Y(N460) );
  NOR3X1TF U439 ( .A(N1056), .B(N1055), .C(N1054), .Y(N1057) );
  OAI22X1TF U440 ( .A0(N642), .A1(N1179), .B0(N674), .B1(N221), .Y(N1055) );
  OAI22X1TF U441 ( .A0(N690), .A1(N1176), .B0(N180), .B1(N1129), .Y(N1056) );
  OAI21X1TF U442 ( .A0(N628), .A1(N148), .B0(N1134), .Y(N496) );
  NOR3X1TF U443 ( .A(N1133), .B(N1132), .C(N1131), .Y(N1134) );
  OAI22X1TF U444 ( .A0(N660), .A1(N222), .B0(N1130), .B1(N1180), .Y(N1131) );
  OAI22X1TF U445 ( .A0(N644), .A1(N1179), .B0(N676), .B1(N221), .Y(N1132) );
  OAI22X1TF U446 ( .A0(N692), .A1(N1176), .B0(N198), .B1(N1129), .Y(N1133) );
  OAI21X1TF U447 ( .A0(N623), .A1(N148), .B0(N920), .Y(N443) );
  NOR3X1TF U448 ( .A(N919), .B(N918), .C(N917), .Y(N920) );
  OAI22X1TF U449 ( .A0(N639), .A1(N1680), .B0(N671), .B1(N221), .Y(N918) );
  OAI22X1TF U450 ( .A0(N687), .A1(N155), .B0(N402), .B1(N1177), .Y(N919) );
  OAI21X1TF U451 ( .A0(N622), .A1(N148), .B0(N916), .Y(N442) );
  NOR3X1TF U452 ( .A(N915), .B(N914), .C(N913), .Y(N916) );
  OAI22X1TF U453 ( .A0(N638), .A1(N1680), .B0(N670), .B1(N221), .Y(N914) );
  OAI22X1TF U454 ( .A0(N686), .A1(N155), .B0(N403), .B1(N1177), .Y(N915) );
  OAI21X1TF U455 ( .A0(N625), .A1(N148), .B0(N1091), .Y(N4780) );
  NOR3X1TF U456 ( .A(N1090), .B(N1089), .C(N1088), .Y(N1091) );
  OAI22X1TF U457 ( .A0(N641), .A1(N1680), .B0(N673), .B1(N221), .Y(N1089) );
  OAI22X1TF U458 ( .A0(N689), .A1(N1176), .B0(N400), .B1(N1129), .Y(N1090) );
  OAI21X1TF U459 ( .A0(N621), .A1(N148), .B0(N1185), .Y(N5140) );
  NOR3X1TF U460 ( .A(N1184), .B(N1183), .C(N1182), .Y(N1185) );
  OAI22X1TF U461 ( .A0(N653), .A1(N222), .B0(N405), .B1(N1180), .Y(N1182) );
  OAI22X1TF U462 ( .A0(N637), .A1(N1680), .B0(N669), .B1(N221), .Y(N1183) );
  OAI22X1TF U463 ( .A0(N404), .A1(N1177), .B0(N685), .B1(N1176), .Y(N1184) );
  OAI21X1TF U464 ( .A0(N420), .A1(N35), .B0(N907), .Y(N440) );
  NOR3X1TF U465 ( .A(N906), .B(N905), .C(N904), .Y(N907) );
  OAI22X1TF U466 ( .A0(N620), .A1(N147), .B0(N652), .B1(N222), .Y(N904) );
  OAI22X1TF U467 ( .A0(N684), .A1(N1176), .B0(N198), .B1(N1152), .Y(N906) );
  OAI21X1TF U468 ( .A0(N418), .A1(N1180), .B0(N899), .Y(N438) );
  NOR3X1TF U469 ( .A(N898), .B(N897), .C(N896), .Y(N899) );
  OAI22X1TF U470 ( .A0(N619), .A1(N147), .B0(N651), .B1(N222), .Y(N896) );
  OAI22X1TF U471 ( .A0(N683), .A1(N1176), .B0(N185), .B1(N1152), .Y(N898) );
  OAI21X1TF U472 ( .A0(N412), .A1(N35), .B0(N891), .Y(N436) );
  NOR3X1TF U473 ( .A(N890), .B(N889), .C(N888), .Y(N891) );
  OAI22X1TF U474 ( .A0(N613), .A1(N147), .B0(N645), .B1(N222), .Y(N888) );
  OAI22X1TF U475 ( .A0(N677), .A1(N1176), .B0(N404), .B1(N1152), .Y(N890) );
  OAI21X1TF U476 ( .A0(N411), .A1(N35), .B0(N1145), .Y(N501) );
  NOR3X1TF U477 ( .A(N1144), .B(N1143), .C(N1142), .Y(N1145) );
  OAI22X1TF U478 ( .A0(N6160), .A1(N147), .B0(N648), .B1(N222), .Y(N1142) );
  OAI22X1TF U479 ( .A0(N632), .A1(N1179), .B0(N664), .B1(N221), .Y(N1143) );
  OAI22X1TF U480 ( .A0(N680), .A1(N1176), .B0(N401), .B1(N1152), .Y(N1144) );
  OAI21X1TF U481 ( .A0(N415), .A1(N35), .B0(N895), .Y(N437) );
  NOR3X1TF U482 ( .A(N894), .B(N893), .C(N892), .Y(N895) );
  OAI22X1TF U483 ( .A0(N614), .A1(N147), .B0(N646), .B1(N222), .Y(N892) );
  OAI22X1TF U484 ( .A0(N678), .A1(N155), .B0(N403), .B1(N1152), .Y(N894) );
  OAI21X1TF U485 ( .A0(N413), .A1(N35), .B0(N903), .Y(N439) );
  NOR3X1TF U486 ( .A(N902), .B(N901), .C(N900), .Y(N903) );
  OAI22X1TF U487 ( .A0(N615), .A1(N147), .B0(N647), .B1(N222), .Y(N900) );
  OAI22X1TF U488 ( .A0(N679), .A1(N155), .B0(N402), .B1(N1152), .Y(N902) );
  OAI21X1TF U489 ( .A0(N408), .A1(N35), .B0(N1081), .Y(N4730) );
  NOR3X1TF U490 ( .A(N1080), .B(N1079), .C(N1078), .Y(N1081) );
  OAI22X1TF U491 ( .A0(N618), .A1(N147), .B0(N650), .B1(N222), .Y(N1078) );
  OAI22X1TF U492 ( .A0(N634), .A1(N1680), .B0(N666), .B1(N221), .Y(N1079) );
  OAI22X1TF U493 ( .A0(N682), .A1(N155), .B0(N180), .B1(N1152), .Y(N1080) );
  OAI21X1TF U494 ( .A0(N409), .A1(N35), .B0(N1156), .Y(N5060) );
  NOR3X1TF U495 ( .A(N1155), .B(N1154), .C(N1153), .Y(N1156) );
  OAI22X1TF U496 ( .A0(N617), .A1(N147), .B0(N649), .B1(N222), .Y(N1153) );
  NOR2X1TF U497 ( .A(OPER3_R3[0]), .B(N886), .Y(N887) );
  OAI22X1TF U498 ( .A0(N633), .A1(N1680), .B0(N665), .B1(N221), .Y(N1154) );
  NOR2X1TF U499 ( .A(OPER3_R3[1]), .B(N886), .Y(N884) );
  INVX2TF U500 ( .A(N885), .Y(N886) );
  OAI22X1TF U501 ( .A0(N681), .A1(N155), .B0(N400), .B1(N1152), .Y(N1155) );
  NAND2X2TF U502 ( .A(N882), .B(N1012), .Y(N1152) );
  AOI211X1TF U503 ( .A0(N729), .A1(N728), .B0(CODE_TYPE[2]), .C0(N1031), .Y(
        N882) );
  OAI211X1TF U504 ( .A0(N880), .A1(N182), .B0(N879), .C0(N878), .Y(N908) );
  INVX2TF U505 ( .A(N1009), .Y(N392) );
  AOI21X1TF U506 ( .A0(N877), .A1(N876), .B0(N875), .Y(N881) );
  AOI21X1TF U507 ( .A0(D_ADDR[2]), .A1(N709), .B0(N612), .Y(N812) );
  OAI21X1TF U508 ( .A0(N703), .A1(N208), .B0(N611), .Y(N612) );
  OAI211X1TF U509 ( .A0(I_ADDR[1]), .A1(I_ADDR[2]), .B0(N700), .C0(N693), .Y(
        N611) );
  AOI211X1TF U510 ( .A0(N709), .A1(D_ADDR[3]), .B0(N695), .C0(N694), .Y(N811)
         );
  AOI211X1TF U511 ( .A0(N693), .A1(N184), .B0(N696), .C0(N704), .Y(N694) );
  NOR2X1TF U512 ( .A(N184), .B(N703), .Y(N695) );
  AOI21X1TF U513 ( .A0(D_ADDR[1]), .A1(N709), .B0(N5190), .Y(N860) );
  AOI22X1TF U514 ( .A0(I_ADDR[1]), .A1(N703), .B0(N704), .B1(N196), .Y(N5190)
         );
  AOI211X1TF U515 ( .A0(N709), .A1(D_ADDR[5]), .B0(N699), .C0(N698), .Y(N809)
         );
  AOI211X1TF U516 ( .A0(N697), .A1(N209), .B0(N701), .C0(N704), .Y(N698) );
  NOR2X1TF U517 ( .A(N209), .B(N703), .Y(N699) );
  AOI211X1TF U518 ( .A0(N709), .A1(D_ADDR[7]), .B0(N708), .C0(N707), .Y(N804)
         );
  AOI211X1TF U519 ( .A0(N706), .A1(N212), .B0(N705), .C0(N704), .Y(N707) );
  NOR2X1TF U520 ( .A(N212), .B(N703), .Y(N708) );
  OAI32X1TF U521 ( .A0(N536), .A1(N705), .A2(I_ADDR[8]), .B0(N700), .B1(N536), 
        .Y(N859) );
  INVX2TF U522 ( .A(N704), .Y(N700) );
  INVX2TF U523 ( .A(N703), .Y(N702) );
  NOR2X1TF U524 ( .A(N697), .B(N209), .Y(N701) );
  NOR3X1TF U525 ( .A(N196), .B(N208), .C(N184), .Y(N696) );
  NOR2X2TF U526 ( .A(N544), .B(N5170), .Y(N709) );
  AOI32X1TF U527 ( .A0(N5150), .A1(N1006), .A2(N211), .B0(N5120), .B1(N1006), 
        .Y(N5170) );
  OAI22X1TF U528 ( .A0(N728), .A1(N211), .B0(N5090), .B1(N5040), .Y(N5120) );
  OAI22X1TF U529 ( .A0(CF), .A1(N877), .B0(N499), .B1(N181), .Y(N5040) );
  AOI21X1TF U530 ( .A0(CF), .A1(N186), .B0(N135), .Y(N499) );
  AOI22X1TF U531 ( .A0(I_ADDR[0]), .A1(N595), .B0(N603), .B1(N193), .Y(
        D_DATAOUT[7]) );
  AOI22X1TF U532 ( .A0(I_ADDR[0]), .A1(N596), .B0(N604), .B1(N193), .Y(
        D_DATAOUT[6]) );
  AOI22X1TF U533 ( .A0(I_ADDR[0]), .A1(N597), .B0(N605), .B1(N193), .Y(
        D_DATAOUT[5]) );
  AOI22X1TF U534 ( .A0(I_ADDR[0]), .A1(N598), .B0(N606), .B1(N193), .Y(
        D_DATAOUT[4]) );
  AOI22X1TF U535 ( .A0(I_ADDR[0]), .A1(N599), .B0(N607), .B1(N193), .Y(
        D_DATAOUT[3]) );
  AOI22X1TF U536 ( .A0(I_ADDR[0]), .A1(N600), .B0(N608), .B1(N193), .Y(
        D_DATAOUT[2]) );
  AOI22X1TF U537 ( .A0(I_ADDR[0]), .A1(N601), .B0(N609), .B1(N193), .Y(
        D_DATAOUT[1]) );
  AOI22X1TF U538 ( .A0(I_ADDR[0]), .A1(N602), .B0(N610), .B1(N193), .Y(
        D_DATAOUT[0]) );
  AOI22X1TF U539 ( .A0(N151), .A1(N1192), .B0(N569), .B1(N1191), .Y(N532) );
  AOI22X1TF U540 ( .A0(N151), .A1(N1190), .B0(N182), .B1(N1191), .Y(N528) );
  AOI22X1TF U541 ( .A0(N149), .A1(N1190), .B0(N404), .B1(N1188), .Y(N520) );
  INVX2TF U542 ( .A(I_DATAIN[7]), .Y(N1190) );
  AOI22X1TF U543 ( .A0(N149), .A1(N1192), .B0(N400), .B1(N1188), .Y(N524) );
  INVX2TF U544 ( .A(I_DATAIN[3]), .Y(N1192) );
  AOI22X1TF U545 ( .A0(N585), .A1(N584), .B0(N629), .B1(N583), .Y(N929) );
  AOI22X1TF U546 ( .A0(N579), .A1(N584), .B0(N661), .B1(N578), .Y(N945) );
  AOI22X1TF U547 ( .A0(N581), .A1(N591), .B0(N647), .B1(N580), .Y(N939) );
  AOI22X1TF U548 ( .A0(N585), .A1(N591), .B0(N631), .B1(N583), .Y(N931) );
  AOI22X1TF U549 ( .A0(N581), .A1(N593), .B0(N646), .B1(N580), .Y(N938) );
  AOI22X1TF U550 ( .A0(N579), .A1(N593), .B0(N662), .B1(N578), .Y(N946) );
  AOI22X1TF U551 ( .A0(N581), .A1(N584), .B0(N645), .B1(N580), .Y(N937) );
  AOI22X1TF U552 ( .A0(N585), .A1(N593), .B0(N630), .B1(N583), .Y(N930) );
  AOI22X1TF U553 ( .A0(N579), .A1(N591), .B0(N663), .B1(N578), .Y(N947) );
  AOI22X1TF U554 ( .A0(N594), .A1(N593), .B0(N614), .B1(N592), .Y(N922) );
  AOI22X1TF U555 ( .A0(N594), .A1(N584), .B0(N613), .B1(N592), .Y(N1001) );
  AOI22X1TF U556 ( .A0(N594), .A1(N591), .B0(N615), .B1(N592), .Y(N923) );
  AOI22X1TF U557 ( .A0(N575), .A1(N591), .B0(N679), .B1(N574), .Y(N955) );
  AOI22X1TF U558 ( .A0(N575), .A1(N593), .B0(N678), .B1(N574), .Y(N954) );
  AOI22X1TF U559 ( .A0(N575), .A1(N584), .B0(N677), .B1(N574), .Y(N953) );
  AOI22X1TF U560 ( .A0(N585), .A1(N590), .B0(N632), .B1(N583), .Y(N932) );
  AOI22X1TF U561 ( .A0(N556), .A1(N562), .B0(N640), .B1(N555), .Y(N972) );
  AOI22X1TF U562 ( .A0(N556), .A1(N563), .B0(N639), .B1(N555), .Y(N971) );
  AOI22X1TF U563 ( .A0(N550), .A1(N558), .B0(N676), .B1(N549), .Y(N992) );
  AOI22X1TF U564 ( .A0(N550), .A1(N563), .B0(N671), .B1(N549), .Y(N987) );
  AOI22X1TF U565 ( .A0(N556), .A1(N558), .B0(N644), .B1(N555), .Y(N976) );
  AOI22X1TF U566 ( .A0(N579), .A1(N5880), .B0(N666), .B1(N578), .Y(N950) );
  AOI22X1TF U567 ( .A0(N579), .A1(N590), .B0(N664), .B1(N578), .Y(N948) );
  AOI22X1TF U568 ( .A0(N550), .A1(N562), .B0(N672), .B1(N549), .Y(N988) );
  AOI22X1TF U569 ( .A0(N550), .A1(N561), .B0(N673), .B1(N549), .Y(N989) );
  AOI22X1TF U570 ( .A0(N550), .A1(N560), .B0(N674), .B1(N549), .Y(N990) );
  INVX2TF U571 ( .A(N550), .Y(N549) );
  AOI22X1TF U572 ( .A0(N581), .A1(N590), .B0(N648), .B1(N580), .Y(N940) );
  AOI22X1TF U573 ( .A0(N556), .A1(N561), .B0(N641), .B1(N555), .Y(N973) );
  AOI22X1TF U574 ( .A0(N594), .A1(N5880), .B0(N618), .B1(N592), .Y(N926) );
  AOI22X1TF U575 ( .A0(N594), .A1(N5890), .B0(N617), .B1(N592), .Y(N925) );
  AOI22X1TF U576 ( .A0(N594), .A1(N590), .B0(N6160), .B1(N592), .Y(N924) );
  AOI22X1TF U577 ( .A0(N594), .A1(N586), .B0(N620), .B1(N592), .Y(N928) );
  AOI22X1TF U578 ( .A0(N594), .A1(N587), .B0(N619), .B1(N592), .Y(N927) );
  NAND4X2TF U579 ( .A(N572), .B(N571), .C(\OPER1_R1[2] ), .D(N576), .Y(N592)
         );
  AOI22X1TF U580 ( .A0(N575), .A1(N590), .B0(N680), .B1(N574), .Y(N956) );
  AOI22X1TF U581 ( .A0(N575), .A1(N5880), .B0(N682), .B1(N574), .Y(N958) );
  AOI22X1TF U582 ( .A0(N575), .A1(N586), .B0(N684), .B1(N574), .Y(N960) );
  AOI22X1TF U583 ( .A0(N575), .A1(N587), .B0(N683), .B1(N574), .Y(N959) );
  AOI22X1TF U584 ( .A0(N575), .A1(N5890), .B0(N681), .B1(N574), .Y(N957) );
  INVX2TF U585 ( .A(N146), .Y(N568) );
  INVX2TF U586 ( .A(N574), .Y(N575) );
  NAND2X2TF U587 ( .A(N576), .B(N1010), .Y(N574) );
  AOI22X1TF U588 ( .A0(N548), .A1(N563), .B0(N687), .B1(N547), .Y(N995) );
  AOI22X1TF U589 ( .A0(N548), .A1(N562), .B0(N688), .B1(N547), .Y(N996) );
  AOI22X1TF U590 ( .A0(N548), .A1(N566), .B0(N685), .B1(N547), .Y(N993) );
  AOI22X1TF U591 ( .A0(N548), .A1(N559), .B0(N691), .B1(N547), .Y(N999) );
  AOI22X1TF U592 ( .A0(N548), .A1(N560), .B0(N690), .B1(N547), .Y(N998) );
  AOI22X1TF U593 ( .A0(N548), .A1(N561), .B0(N689), .B1(N547), .Y(N997) );
  AOI22X1TF U594 ( .A0(N548), .A1(N558), .B0(N692), .B1(N547), .Y(N1000) );
  AOI22X1TF U595 ( .A0(N548), .A1(N564), .B0(N686), .B1(N547), .Y(N994) );
  AOI22X1TF U596 ( .A0(N552), .A1(N563), .B0(N655), .B1(N551), .Y(N979) );
  AOI22X1TF U597 ( .A0(N552), .A1(N558), .B0(N660), .B1(N551), .Y(N984) );
  AOI22X1TF U598 ( .A0(N552), .A1(N562), .B0(N656), .B1(N551), .Y(N980) );
  AOI22X1TF U599 ( .A0(N552), .A1(N566), .B0(N653), .B1(N551), .Y(N977) );
  AOI22X1TF U600 ( .A0(N552), .A1(N561), .B0(N657), .B1(N551), .Y(N981) );
  AOI22X1TF U601 ( .A0(N552), .A1(N564), .B0(N654), .B1(N551), .Y(N978) );
  AOI22X1TF U602 ( .A0(N567), .A1(N558), .B0(N628), .B1(N565), .Y(N968) );
  AOI22X1TF U603 ( .A0(N567), .A1(N563), .B0(N623), .B1(N565), .Y(N963) );
  AOI22X1TF U604 ( .A0(N567), .A1(N562), .B0(N624), .B1(N565), .Y(N964) );
  AOI22X1TF U605 ( .A0(N567), .A1(N561), .B0(N625), .B1(N565), .Y(N965) );
  AOI22X1TF U606 ( .A0(N567), .A1(N564), .B0(N622), .B1(N565), .Y(N962) );
  AOI22X1TF U607 ( .A0(N567), .A1(N566), .B0(N621), .B1(N565), .Y(N961) );
  AOI22X1TF U608 ( .A0(N567), .A1(N559), .B0(N627), .B1(N565), .Y(N967) );
  AOI22X1TF U609 ( .A0(N567), .A1(N560), .B0(N626), .B1(N565), .Y(N966) );
  NAND4X2TF U610 ( .A(N571), .B(N572), .C(\OPER1_R1[2] ), .D(N557), .Y(N565)
         );
  INVX2TF U611 ( .A(N573), .Y(N543) );
  NOR2X1TF U612 ( .A(N217), .B(N545), .Y(N537) );
  OAI211X1TF U613 ( .A0(STATE[1]), .A1(N721), .B0(I_ADDR[0]), .C0(N873), .Y(
        N538) );
  INVX2TF U614 ( .A(N712), .Y(N721) );
  AOI21X1TF U615 ( .A0(N357), .A1(N1173), .B0(N355), .Y(N356) );
  OAI21X1TF U616 ( .A0(N374), .A1(N125), .B0(N354), .Y(N355) );
  AOI22X1TF U617 ( .A0(IO_DATAINB[8]), .A1(N220), .B0(REG_C[8]), .B1(N1172), 
        .Y(N354) );
  AOI21X1TF U618 ( .A0(N352), .A1(N1175), .B0(N351), .Y(N353) );
  AOI22X1TF U619 ( .A0(IO_DATAINB[4]), .A1(N220), .B0(D_ADDR[5]), .B1(N1172), 
        .Y(N349) );
  OAI211X1TF U620 ( .A0(N361), .A1(N127), .B0(N359), .C0(N358), .Y(N360) );
  AOI21X1TF U621 ( .A0(N512), .A1(N218), .B0(N335), .Y(N336) );
  OAI21X1TF U622 ( .A0(N826), .A1(N816), .B0(N334), .Y(N335) );
  OAI22X1TF U623 ( .A0(N829), .A1(N831), .B0(N819), .B1(N869), .Y(N332) );
  OAI22X1TF U624 ( .A0(N820), .A1(N828), .B0(N827), .B1(N862), .Y(N818) );
  NOR2X1TF U625 ( .A(N331), .B(N206), .Y(N333) );
  AOI22X1TF U626 ( .A0(REG_A[8]), .A1(N390), .B0(N389), .B1(N206), .Y(N814) );
  AOI22X1TF U627 ( .A0(IO_DATAINB[9]), .A1(N220), .B0(REG_C[9]), .B1(N1172), 
        .Y(N359) );
  AOI22X1TF U628 ( .A0(N1141), .A1(IO_STATUS[1]), .B0(N169), .B1(IO_DATAINA[1]), .Y(N1121) );
  AOI22X1TF U629 ( .A0(IO_DATAINB[1]), .A1(N378), .B0(D_ADDR[2]), .B1(N150), 
        .Y(N1122) );
  AOI21X1TF U630 ( .A0(N479), .A1(N219), .B0(N288), .Y(N361) );
  AOI211X1TF U631 ( .A0(REG_A[9]), .A1(N286), .B0(N802), .C0(N285), .Y(N287)
         );
  OAI21X1TF U632 ( .A0(N800), .A1(N826), .B0(N284), .Y(N285) );
  AOI211X1TF U633 ( .A0(N852), .A1(N837), .B0(N283), .C0(N803), .Y(N284) );
  OAI22X1TF U634 ( .A0(N835), .A1(N828), .B0(N798), .B1(N203), .Y(N803) );
  NOR2X1TF U635 ( .A(N862), .B(N801), .Y(N283) );
  AOI22X1TF U636 ( .A0(REG_A[9]), .A1(N152), .B0(N225), .B1(N176), .Y(N799) );
  AOI21X1TF U637 ( .A0(N481), .A1(N219), .B0(N276), .Y(N372) );
  AOI211X1TF U638 ( .A0(REG_A[11]), .A1(N274), .B0(N273), .C0(N754), .Y(N275)
         );
  AOI22X1TF U639 ( .A0(REG_A[11]), .A1(N390), .B0(N225), .B1(N194), .Y(N751)
         );
  OAI21X1TF U640 ( .A0(N753), .A1(N862), .B0(N272), .Y(N273) );
  AOI211X1TF U641 ( .A0(N752), .A1(N325), .B0(N271), .C0(N755), .Y(N272) );
  OAI22X1TF U642 ( .A0(N789), .A1(N869), .B0(N828), .B1(N792), .Y(N755) );
  NOR2X1TF U643 ( .A(N831), .B(N797), .Y(N271) );
  OAI211X1TF U644 ( .A0(N380), .A1(N126), .B0(N11000), .C0(N1099), .Y(N4820)
         );
  AOI22X1TF U645 ( .A0(IO_DATAINA[3]), .A1(N169), .B0(N1173), .B1(N352), .Y(
        N1099) );
  OAI211X1TF U646 ( .A0(N797), .A1(N834), .B0(N796), .C0(N341), .Y(N352) );
  OAI21X1TF U647 ( .A0(N789), .A1(N826), .B0(N339), .Y(N340) );
  AOI21X1TF U648 ( .A0(N507), .A1(N863), .B0(N338), .Y(N339) );
  AOI211X1TF U649 ( .A0(REG_A[5]), .A1(N26), .B0(N786), .C0(N785), .Y(N788) );
  AOI221X1TF U650 ( .A0(N1092), .A1(N389), .B0(REG_A[3]), .B1(N152), .C0(N793), 
        .Y(N794) );
  OAI21X1TF U651 ( .A0(REG_B[3]), .A1(N121), .B0(N791), .Y(N795) );
  AOI22X1TF U652 ( .A0(IO_DATAINB[3]), .A1(N378), .B0(D_ADDR[4]), .B1(N1172), 
        .Y(N11000) );
  AOI21X1TF U653 ( .A0(N376), .A1(N1175), .B0(N375), .Y(N377) );
  OAI21X1TF U654 ( .A0(N374), .A1(N127), .B0(N373), .Y(N375) );
  AOI22X1TF U655 ( .A0(IO_DATAINB[7]), .A1(N378), .B0(D_ADDR[8]), .B1(N1172), 
        .Y(N373) );
  AOI21X1TF U656 ( .A0(N477), .A1(N337), .B0(N313), .Y(N374) );
  AOI211X1TF U657 ( .A0(REG_A[7]), .A1(N311), .B0(N749), .C0(N310), .Y(N312)
         );
  OAI211X1TF U658 ( .A0(N797), .A1(N828), .B0(N309), .C0(N308), .Y(N310) );
  OAI22X1TF U659 ( .A0(N789), .A1(N862), .B0(N792), .B1(N834), .Y(N750) );
  INVX2TF U660 ( .A(N740), .Y(N789) );
  NOR4BX1TF U661 ( .AN(N744), .B(N743), .C(N742), .D(N741), .Y(N790) );
  AOI211X1TF U662 ( .A0(REG_A[11]), .A1(N393), .B0(N748), .C0(N747), .Y(N797)
         );
  OAI22X1TF U663 ( .A0(N768), .A1(N1101), .B0(N851), .B1(N178), .Y(N747) );
  INVX2TF U664 ( .A(N746), .Y(N748) );
  AOI22X1TF U665 ( .A0(REG_A[7]), .A1(N152), .B0(N225), .B1(N189), .Y(N745) );
  OAI211X1TF U666 ( .A0(N379), .A1(N128), .B0(N1034), .C0(N1033), .Y(N447) );
  AOI22X1TF U667 ( .A0(IO_DATAINA[5]), .A1(N169), .B0(N1175), .B1(N350), .Y(
        N1033) );
  OR2X2TF U668 ( .A(N830), .B(N330), .Y(N350) );
  AOI22X1TF U669 ( .A0(N474), .A1(N337), .B0(N863), .B1(N508), .Y(N323) );
  OAI22X1TF U670 ( .A0(N820), .A1(N834), .B0(N862), .B1(N819), .Y(N832) );
  INVX2TF U671 ( .A(N815), .Y(N819) );
  INVX2TF U672 ( .A(N845), .Y(N820) );
  INVX2TF U673 ( .A(N847), .Y(N829) );
  AOI22X1TF U674 ( .A0(REG_A[4]), .A1(N152), .B0(N389), .B1(N202), .Y(N825) );
  AOI22X1TF U675 ( .A0(IO_DATAINB[5]), .A1(N378), .B0(D_ADDR[6]), .B1(N150), 
        .Y(N1034) );
  OAI211X1TF U676 ( .A0(N382), .A1(N126), .B0(N1065), .C0(N1064), .Y(N464) );
  INVX2TF U677 ( .A(N344), .Y(N380) );
  OAI211X1TF U678 ( .A0(N870), .A1(N826), .B0(N782), .C0(N315), .Y(N344) );
  AOI211X1TF U679 ( .A0(N506), .A1(N863), .B0(N783), .C0(N314), .Y(N315) );
  INVX2TF U680 ( .A(N773), .Y(N784) );
  OAI22X1TF U681 ( .A0(N779), .A1(N831), .B0(N865), .B1(N778), .Y(N783) );
  AOI211X1TF U682 ( .A0(REG_A[4]), .A1(N26), .B0(N775), .C0(N774), .Y(N779) );
  AOI22X1TF U683 ( .A0(REG_B[2]), .A1(N781), .B0(REG_A[2]), .B1(N780), .Y(N782) );
  OAI21X1TF U684 ( .A0(REG_B[2]), .A1(N121), .B0(N791), .Y(N780) );
  AOI22X1TF U685 ( .A0(IO_DATAINB[2]), .A1(N378), .B0(D_ADDR[3]), .B1(N150), 
        .Y(N1065) );
  INVX2TF U686 ( .A(N345), .Y(N382) );
  AOI21X1TF U687 ( .A0(N471), .A1(N219), .B0(N317), .Y(N319) );
  OAI211X1TF U688 ( .A0(N202), .A1(N768), .B0(N767), .C0(N766), .Y(N769) );
  OAI32X1TF U689 ( .A0(N1112), .A1(REG_B[1]), .A2(N121), .B0(N791), .B1(N1112), 
        .Y(N771) );
  AOI21X1TF U690 ( .A0(N376), .A1(N1173), .B0(N347), .Y(N348) );
  OAI21X1TF U691 ( .A0(N379), .A1(N126), .B0(N346), .Y(N347) );
  AOI22X1TF U692 ( .A0(IO_DATAINB[6]), .A1(N220), .B0(D_ADDR[7]), .B1(N1172), 
        .Y(N346) );
  AOI211X1TF U693 ( .A0(N475), .A1(N219), .B0(N306), .C0(N305), .Y(N379) );
  AOI211X1TF U694 ( .A0(N839), .A1(N303), .B0(N840), .C0(N302), .Y(N304) );
  OAI22X1TF U695 ( .A0(N835), .A1(N834), .B0(N833), .B1(N836), .Y(N840) );
  OAI21X1TF U696 ( .A0(N826), .A1(N861), .B0(N294), .Y(N376) );
  AOI211X1TF U697 ( .A0(N476), .A1(N337), .B0(N293), .C0(N738), .Y(N294) );
  AOI22X1TF U698 ( .A0(REG_A[6]), .A1(N152), .B0(N225), .B1(N207), .Y(N734) );
  OAI211X1TF U699 ( .A0(N292), .A1(N207), .B0(N291), .C0(N290), .Y(N293) );
  AOI211X1TF U700 ( .A0(N838), .A1(N776), .B0(N289), .C0(N739), .Y(N290) );
  OAI22X1TF U701 ( .A0(N870), .A1(N862), .B0(N730), .B1(N778), .Y(N739) );
  NOR2X1TF U702 ( .A(N831), .B(N773), .Y(N289) );
  INVX2TF U703 ( .A(N828), .Y(N838) );
  AOI21X1TF U704 ( .A0(IO_DATAINA[0]), .A1(N169), .B0(N368), .Y(N369) );
  OAI211X1TF U705 ( .A0(N381), .A1(N127), .B0(N367), .C0(N366), .Y(N368) );
  NOR2X1TF U706 ( .A(N24), .B(N1119), .Y(N1141) );
  AOI22X1TF U707 ( .A0(IO_DATAINB[0]), .A1(N220), .B0(D_ADDR[1]), .B1(N1172), 
        .Y(N367) );
  AND2X2TF U708 ( .A(N217), .B(N343), .Y(N378) );
  AND2X2TF U709 ( .A(N391), .B(N342), .Y(N343) );
  INVX2TF U710 ( .A(N1030), .Y(N342) );
  AOI211X1TF U711 ( .A0(REG_A[0]), .A1(N300), .B0(N299), .C0(N298), .Y(N381)
         );
  OAI211X1TF U712 ( .A0(N857), .A1(N858), .B0(N856), .C0(N297), .Y(N298) );
  AOI22X1TF U713 ( .A0(N218), .A1(N504), .B0(N470), .B1(N219), .Y(N297) );
  OAI31X1TF U714 ( .A0(N855), .A1(N854), .A2(N853), .B0(N852), .Y(N856) );
  NOR2X1TF U715 ( .A(N851), .B(N177), .Y(N853) );
  NOR2X1TF U716 ( .A(N850), .B(N1112), .Y(N854) );
  OAI22X1TF U717 ( .A0(REG_A[0]), .A1(N121), .B0(N842), .B1(N187), .Y(N296) );
  OAI21X1TF U718 ( .A0(REG_B[0]), .A1(N121), .B0(N295), .Y(N300) );
  OAI211X1TF U719 ( .A0(N861), .A1(N862), .B0(N281), .C0(N280), .Y(N282) );
  NOR3X1TF U720 ( .A(N279), .B(N871), .C(N278), .Y(N280) );
  AOI22X1TF U721 ( .A0(REG_B[2]), .A1(N777), .B0(N776), .B1(N201), .Y(N865) );
  OAI211X1TF U722 ( .A0(N124), .A1(N188), .B0(N737), .C0(N736), .Y(N776) );
  INVX2TF U723 ( .A(N857), .Y(N864) );
  OAI22X1TF U724 ( .A0(N870), .A1(N869), .B0(N868), .B1(N188), .Y(N871) );
  OAI211X1TF U725 ( .A0(N417), .A1(N411), .B0(N256), .C0(N255), .Y(N257) );
  AOI211X1TF U726 ( .A0(REG_A[12]), .A1(N254), .B0(N253), .C0(N252), .Y(N255)
         );
  OAI211X1TF U727 ( .A0(N190), .A1(N124), .B0(N422), .C0(N398), .Y(N845) );
  OAI211X1TF U728 ( .A0(N176), .A1(N768), .B0(N737), .C0(N806), .Y(N397) );
  NOR2X1TF U729 ( .A(N765), .B(N419), .Y(N253) );
  INVX2TF U730 ( .A(N827), .Y(N407) );
  AOI211X1TF U731 ( .A0(REG_A[4]), .A1(N393), .B0(N775), .C0(N399), .Y(N827)
         );
  OAI22X1TF U732 ( .A0(N768), .A1(N1112), .B0(N851), .B1(N177), .Y(N399) );
  NOR2X1TF U733 ( .A(N850), .B(N1092), .Y(N775) );
  NOR2X1TF U734 ( .A(N124), .B(N187), .Y(N815) );
  INVX2TF U735 ( .A(N816), .Y(N410) );
  NOR4X1TF U736 ( .A(N731), .B(N774), .C(N813), .D(N822), .Y(N816) );
  NOR2X1TF U737 ( .A(N207), .B(N851), .Y(N822) );
  NOR2X1TF U738 ( .A(N123), .B(N206), .Y(N813) );
  NOR2X1TF U739 ( .A(N768), .B(N836), .Y(N774) );
  NOR2X1TF U740 ( .A(N850), .B(N189), .Y(N731) );
  INVX2TF U741 ( .A(N121), .Y(N225) );
  AOI211X1TF U742 ( .A0(REG_A[13]), .A1(N248), .B0(N247), .C0(N246), .Y(N249)
         );
  OAI21X1TF U743 ( .A0(N835), .A1(N831), .B0(N245), .Y(N246) );
  AOI211X1TF U744 ( .A0(N244), .A1(N839), .B0(N243), .C0(N242), .Y(N245) );
  AOI31X1TF U745 ( .A0(N760), .A1(N746), .A2(N744), .B0(N826), .Y(N242) );
  NOR2X1TF U746 ( .A(N862), .B(N800), .Y(N243) );
  NOR4BBX1TF U747 ( .AN(N756), .BN(N761), .C(N741), .D(N785), .Y(N800) );
  NOR2X1TF U748 ( .A(N207), .B(N768), .Y(N785) );
  NOR2X1TF U749 ( .A(N206), .B(N850), .Y(N741) );
  OAI22X1TF U750 ( .A0(N201), .A1(N764), .B0(N801), .B1(REG_B[2]), .Y(N839) );
  AOI211X1TF U751 ( .A0(REG_A[2]), .A1(N735), .B0(N394), .C0(N786), .Y(N801)
         );
  NOR2X1TF U752 ( .A(N850), .B(N202), .Y(N786) );
  OAI22X1TF U753 ( .A0(N124), .A1(N836), .B0(N851), .B1(N1092), .Y(N394) );
  INVX2TF U754 ( .A(N798), .Y(N244) );
  AOI21X1TF U755 ( .A0(N393), .A1(REG_A[13]), .B0(N395), .Y(N835) );
  OAI22X1TF U756 ( .A0(N851), .A1(N192), .B0(N850), .B1(N1101), .Y(N395) );
  NOR3X1TF U757 ( .A(N730), .B(REG_B[3]), .C(N857), .Y(N258) );
  AOI221X1TF U758 ( .A0(REG_B[0]), .A1(N192), .B0(N1130), .B1(N1101), .C0(
        REG_B[1]), .Y(N777) );
  AOI31X1TF U759 ( .A0(N425), .A1(N805), .A2(N422), .B0(N826), .Y(N450) );
  OAI22X1TF U760 ( .A0(N432), .A1(N765), .B0(N415), .B1(N431), .Y(N446) );
  INVX2TF U761 ( .A(N870), .Y(N429) );
  AOI21X1TF U762 ( .A0(N393), .A1(REG_A[2]), .B0(N428), .Y(N870) );
  OAI22X1TF U763 ( .A0(N851), .A1(N187), .B0(N850), .B1(N1112), .Y(N428) );
  NOR4X1TF U764 ( .A(N732), .B(N855), .C(N426), .D(N823), .Y(N861) );
  NOR2X1TF U765 ( .A(N850), .B(N836), .Y(N823) );
  INVX2TF U766 ( .A(N467), .Y(N850) );
  NOR2X1TF U767 ( .A(N851), .B(N202), .Y(N426) );
  NOR2X1TF U768 ( .A(N768), .B(N1092), .Y(N855) );
  NOR2X1TF U769 ( .A(N207), .B(N123), .Y(N732) );
  AOI32X1TF U770 ( .A0(N389), .A1(REG_A[14]), .A2(N415), .B0(N458), .B1(
        REG_A[14]), .Y(N454) );
  INVX2TF U771 ( .A(N396), .Y(N251) );
  OAI21X1TF U772 ( .A0(N269), .A1(N192), .B0(N268), .Y(N270) );
  AOI211X1TF U773 ( .A0(N267), .A1(N752), .B0(N266), .C0(N265), .Y(N268) );
  AOI21X1TF U774 ( .A0(N264), .A1(N263), .B0(N826), .Y(N265) );
  AOI22X1TF U775 ( .A0(REG_A[14]), .A1(N467), .B0(REG_A[13]), .B1(N26), .Y(
        N264) );
  NOR2X1TF U776 ( .A(N262), .B(N765), .Y(N266) );
  INVX2TF U777 ( .A(N387), .Y(N765) );
  NOR2X1TF U778 ( .A(N204), .B(N201), .Y(N844) );
  OAI211X1TF U779 ( .A0(N1092), .A1(N124), .B0(N767), .C0(N463), .Y(N740) );
  NOR2X2TF U780 ( .A(REG_B[2]), .B(N204), .Y(N846) );
  INVX2TF U781 ( .A(N753), .Y(N307) );
  NOR4BX1TF U782 ( .AN(N759), .B(N743), .C(N4760), .D(N4710), .Y(N753) );
  NOR2X1TF U783 ( .A(N851), .B(N836), .Y(N4710) );
  NOR2X1TF U784 ( .A(N768), .B(N202), .Y(N4760) );
  INVX2TF U785 ( .A(N735), .Y(N768) );
  NOR2X1TF U786 ( .A(N124), .B(N189), .Y(N743) );
  NOR2X2TF U787 ( .A(N1130), .B(REG_B[1]), .Y(N467) );
  NOR2X1TF U788 ( .A(N176), .B(N851), .Y(N742) );
  INVX2TF U789 ( .A(N787), .Y(N851) );
  INVX2TF U790 ( .A(N862), .Y(N267) );
  NAND2X2TF U791 ( .A(N387), .B(N848), .Y(N862) );
  AOI21X1TF U792 ( .A0(N412), .A1(N224), .B0(N261), .Y(N269) );
  INVX2TF U793 ( .A(N295), .Y(N261) );
  INVX2TF U794 ( .A(N852), .Y(N831) );
  INVX2TF U795 ( .A(N826), .Y(N325) );
  OR2X2TF U796 ( .A(N316), .B(REG_B[2]), .Y(N826) );
  AND2X2TF U797 ( .A(N1032), .B(N229), .Y(N387) );
  AND2X2TF U798 ( .A(N135), .B(N921), .Y(N229) );
  INVX2TF U799 ( .A(N874), .Y(N1030) );
  INVX2TF U800 ( .A(N121), .Y(N224) );
  OAI211X1TF U801 ( .A0(N880), .A1(N1031), .B0(N867), .C0(N396), .Y(N4850) );
  INVX2TF U802 ( .A(N1032), .Y(N877) );
  NOR3X1TF U803 ( .A(N186), .B(N879), .C(N1005), .Y(N1015) );
  INVX2TF U804 ( .A(N1006), .Y(N879) );
  OR2X2TF U805 ( .A(N233), .B(N232), .Y(N863) );
  NOR2X1TF U806 ( .A(N729), .B(N1031), .Y(N232) );
  INVX2TF U807 ( .A(N391), .Y(N1031) );
  OR2X2TF U808 ( .A(N1009), .B(N24), .Y(N729) );
  AOI21X1TF U809 ( .A0(N231), .A1(N876), .B0(N1004), .Y(N233) );
  INVX2TF U810 ( .A(N1005), .Y(N230) );
  NAND2BX2TF U811 ( .AN(CODE_TYPE[4]), .B(CODE_TYPE[3]), .Y(N1004) );
  AOI211X1TF U812 ( .A0(CODE_TYPE[2]), .A1(N237), .B0(CODE_TYPE[3]), .C0(N236), 
        .Y(N238) );
  INVX2TF U813 ( .A(N1007), .Y(N236) );
  OAI21X1TF U814 ( .A0(N24), .A1(N191), .B0(N234), .Y(N235) );
  INVX2TF U815 ( .A(N5150), .Y(N234) );
  NOR2X1TF U816 ( .A(N569), .B(N223), .Y(N5150) );
  INVX2TF U817 ( .A(N540), .Y(N227) );
  OAI22X1TF U818 ( .A0(N648), .A1(N138), .B0(N136), .B1(N6160), .Y(N1146) );
  OAI22X1TF U819 ( .A0(N664), .A1(N131), .B0(N129), .B1(N190), .Y(N1147) );
  OAI22X1TF U820 ( .A0(N649), .A1(N138), .B0(N137), .B1(N617), .Y(N1157) );
  OAI22X1TF U821 ( .A0(N665), .A1(N131), .B0(N130), .B1(N194), .Y(N1158) );
  OAI22X1TF U822 ( .A0(N645), .A1(N138), .B0(N137), .B1(N613), .Y(N1123) );
  OAI22X1TF U823 ( .A0(N661), .A1(N132), .B0(N130), .B1(N192), .Y(N1124) );
  OAI22X1TF U824 ( .A0(N652), .A1(N138), .B0(N137), .B1(N620), .Y(N1048) );
  OAI22X1TF U825 ( .A0(N668), .A1(N132), .B0(N130), .B1(N206), .Y(N1049) );
  OAI22X1TF U826 ( .A0(N658), .A1(N138), .B0(N137), .B1(N626), .Y(N1058) );
  OAI22X1TF U827 ( .A0(N674), .A1(N131), .B0(N130), .B1(N177), .Y(N1059) );
  OAI22X1TF U828 ( .A0(N650), .A1(N139), .B0(N137), .B1(N618), .Y(N1082) );
  OAI22X1TF U829 ( .A0(N666), .A1(N132), .B0(N130), .B1(N188), .Y(N1083) );
  OAI22X1TF U830 ( .A0(N651), .A1(N139), .B0(N136), .B1(N619), .Y(N1072) );
  OAI22X1TF U831 ( .A0(N667), .A1(N132), .B0(N129), .B1(N176), .Y(N1073) );
  OAI22X1TF U832 ( .A0(N653), .A1(N138), .B0(N136), .B1(N621), .Y(N1168) );
  OAI22X1TF U833 ( .A0(N669), .A1(N132), .B0(N129), .B1(N189), .Y(N1169) );
  OAI22X1TF U834 ( .A0(N647), .A1(N139), .B0(N136), .B1(N615), .Y(N1066) );
  OAI22X1TF U835 ( .A0(N663), .A1(N132), .B0(N129), .B1(N178), .Y(N1067) );
  OAI22X1TF U836 ( .A0(N646), .A1(N139), .B0(N136), .B1(N614), .Y(N1102) );
  OAI22X1TF U837 ( .A0(N662), .A1(N132), .B0(N129), .B1(N1101), .Y(N1103) );
  OAI22X1TF U838 ( .A0(N657), .A1(N139), .B0(N137), .B1(N625), .Y(N1093) );
  OAI22X1TF U839 ( .A0(N673), .A1(N132), .B0(N129), .B1(N1092), .Y(N1094) );
  OAI22X1TF U840 ( .A0(N659), .A1(N138), .B0(N137), .B1(N627), .Y(N1113) );
  OAI22X1TF U841 ( .A0(N675), .A1(N131), .B0(N130), .B1(N1112), .Y(N1114) );
  OAI22X1TF U842 ( .A0(N660), .A1(N138), .B0(N137), .B1(N628), .Y(N1135) );
  OAI22X1TF U843 ( .A0(N676), .A1(N131), .B0(N130), .B1(N187), .Y(N1136) );
  OAI22X1TF U844 ( .A0(N655), .A1(N139), .B0(N136), .B1(N623), .Y(N1024) );
  OAI22X1TF U845 ( .A0(N654), .A1(N139), .B0(N136), .B1(N622), .Y(N1035) );
  OAI22X1TF U846 ( .A0(N656), .A1(N139), .B0(N136), .B1(N624), .Y(N1041) );
  AOI21X1TF U847 ( .A0(N224), .A1(N420), .B0(N122), .Y(N331) );
  AOI21X1TF U848 ( .A0(N133), .A1(N814), .B0(N420), .Y(N817) );
  AOI21X1TF U849 ( .A0(N133), .A1(N799), .B0(N418), .Y(N802) );
  AOI21X1TF U850 ( .A0(N133), .A1(N751), .B0(N409), .Y(N754) );
  OAI31X1TF U851 ( .A0(N201), .A1(N857), .A2(N792), .B0(N134), .Y(N793) );
  AOI21X1TF U852 ( .A0(N134), .A1(N745), .B0(N405), .Y(N749) );
  AOI21X1TF U853 ( .A0(N134), .A1(N825), .B0(N423), .Y(N830) );
  AOI21X1TF U854 ( .A0(N393), .A1(N852), .B0(N122), .Y(N791) );
  AOI21X1TF U855 ( .A0(N225), .A1(N424), .B0(N122), .Y(N833) );
  AOI21X1TF U856 ( .A0(N134), .A1(N301), .B0(N424), .Y(N306) );
  AOI22X1TF U857 ( .A0(N152), .A1(REG_A[5]), .B0(N224), .B1(N836), .Y(N301) );
  AOI21X1TF U858 ( .A0(N134), .A1(N734), .B0(N406), .Y(N738) );
  AOI21X1TF U859 ( .A0(N224), .A1(N406), .B0(N122), .Y(N292) );
  AOI21X1TF U860 ( .A0(N225), .A1(N408), .B0(N122), .Y(N868) );
  AOI21X1TF U861 ( .A0(N133), .A1(N277), .B0(N408), .Y(N279) );
  AOI22X1TF U862 ( .A0(N390), .A1(REG_A[10]), .B0(N224), .B1(N188), .Y(N277)
         );
  AOI22X1TF U863 ( .A0(N735), .A1(REG_A[15]), .B0(N26), .B1(REG_A[14]), .Y(
        N398) );
  AOI221X1TF U864 ( .A0(N152), .A1(REG_A[12]), .B0(N389), .B1(N190), .C0(N25), 
        .Y(N417) );
  AOI21X1TF U865 ( .A0(N134), .A1(N241), .B0(N413), .Y(N247) );
  AOI22X1TF U866 ( .A0(N152), .A1(REG_A[13]), .B0(N224), .B1(N178), .Y(N241)
         );
  AOI221X1TF U867 ( .A0(N152), .A1(REG_A[14]), .B0(N389), .B1(N1101), .C0(N25), 
        .Y(N431) );
  MXI2X1TF U868 ( .A(N362), .B(N211), .S0(N1187), .Y(N435) );
  NAND2X1TF U869 ( .A(OPER3_R3[1]), .B(N887), .Y(N1181) );
  NAND2X1TF U870 ( .A(OPER3_R3[0]), .B(N884), .Y(N1178) );
  OAI32XLTF U871 ( .A0(ZF), .A1(N186), .A2(N876), .B0(N729), .B1(N213), .Y(
        N5090) );
  INVX2TF U872 ( .A(N1016), .Y(N577) );
  INVX2TF U873 ( .A(N547), .Y(N548) );
  OAI2BB1X1TF U874 ( .A0N(N169), .A1N(IO_DATAINA[8]), .B0(N356), .Y(N459) );
  OAI2BB1X1TF U875 ( .A0N(N169), .A1N(IO_DATAINA[4]), .B0(N353), .Y(N455) );
  OAI2BB1X1TF U876 ( .A0N(N1173), .A1N(N350), .B0(N349), .Y(N351) );
  NAND2X1TF U877 ( .A(N357), .B(N1175), .Y(N358) );
  OAI2BB1X1TF U878 ( .A0N(N863), .A1N(N513), .B0(N287), .Y(N288) );
  AO21X1TF U879 ( .A0(N224), .A1(N418), .B0(N122), .Y(N286) );
  OAI2BB1X1TF U880 ( .A0N(N218), .A1N(N515), .B0(N275), .Y(N276) );
  AO21X1TF U881 ( .A0(N224), .A1(N409), .B0(N122), .Y(N274) );
  AOI2BB1X1TF U882 ( .A0N(N828), .A1N(N790), .B0(N340), .Y(N341) );
  OAI2BB2XLTF U883 ( .B0(N788), .B1(N831), .A0N(N473), .A1N(N219), .Y(N338) );
  OAI2BB1X1TF U884 ( .A0N(N169), .A1N(IO_DATAINA[7]), .B0(N377), .Y(N5130) );
  OAI2BB1X1TF U885 ( .A0N(N218), .A1N(N511), .B0(N312), .Y(N313) );
  AOI2BB1X1TF U886 ( .A0N(N790), .A1N(N831), .B0(N750), .Y(N308) );
  NAND2X1TF U887 ( .A(N307), .B(N325), .Y(N309) );
  AO21X1TF U888 ( .A0(N389), .A1(N405), .B0(N122), .Y(N311) );
  NAND4X1TF U889 ( .A(N329), .B(N328), .C(N327), .D(N326), .Y(N330) );
  NAND2BX1TF U890 ( .AN(N843), .B(N852), .Y(N326) );
  NAND2BX1TF U891 ( .AN(N827), .B(N325), .Y(N327) );
  AOI2BB1X1TF U892 ( .A0N(N829), .A1N(N828), .B0(N324), .Y(N328) );
  NAND2BX1TF U893 ( .AN(N832), .B(N323), .Y(N324) );
  NAND2X1TF U894 ( .A(N322), .B(REG_A[4]), .Y(N329) );
  AO21X1TF U895 ( .A0(N389), .A1(N423), .B0(N122), .Y(N322) );
  AO22X1TF U896 ( .A0(N219), .A1(N472), .B0(N784), .B1(N838), .Y(N314) );
  OAI2BB1X1TF U897 ( .A0N(REG_B[1]), .A1N(N772), .B0(N321), .Y(N345) );
  AOI2BB1X1TF U898 ( .A0N(N770), .A1N(N857), .B0(N320), .Y(N321) );
  NAND3BX1TF U899 ( .AN(N771), .B(N319), .C(N318), .Y(N320) );
  NAND2X1TF U900 ( .A(N218), .B(N505), .Y(N318) );
  OAI2BB2XLTF U901 ( .B0(N316), .B1(N203), .A0N(N852), .A1N(N769), .Y(N317) );
  OAI2BB1X1TF U902 ( .A0N(N169), .A1N(IO_DATAINA[6]), .B0(N348), .Y(N451) );
  OAI2BB1X1TF U903 ( .A0N(N509), .A1N(N863), .B0(N304), .Y(N305) );
  AO22X1TF U904 ( .A0(N837), .A1(N838), .B0(N852), .B1(N841), .Y(N302) );
  NAND4X1TF U905 ( .A(N263), .B(N760), .C(N761), .D(N762), .Y(N837) );
  NAND2X1TF U906 ( .A(N510), .B(N863), .Y(N291) );
  NAND2X1TF U907 ( .A(N1141), .B(IO_STATUS[0]), .Y(N366) );
  OA21XLTF U908 ( .A0(N25), .A1(N296), .B0(REG_B[0]), .Y(N299) );
  OAI2BB2XLTF U909 ( .B0(N866), .B1(N865), .A0N(N872), .A1N(N325), .Y(N278) );
  NAND2X1TF U910 ( .A(N514), .B(N218), .Y(N281) );
  AO22X1TF U911 ( .A0(N325), .A1(N397), .B0(N852), .B1(N845), .Y(N252) );
  AOI222XLTF U912 ( .A0(N410), .A1(N848), .B0(N844), .B1(N815), .C0(N407), 
        .C1(N846), .Y(N419) );
  AO21X1TF U913 ( .A0(N225), .A1(N411), .B0(N458), .Y(N254) );
  NAND2X1TF U914 ( .A(N516), .B(N218), .Y(N256) );
  OAI2BB1X1TF U915 ( .A0N(N218), .A1N(N517), .B0(N249), .Y(N250) );
  NAND2X1TF U916 ( .A(N387), .B(REG_B[3]), .Y(N798) );
  AO21X1TF U917 ( .A0(N224), .A1(N413), .B0(N458), .Y(N248) );
  NAND2X1TF U918 ( .A(N735), .B(REG_A[12]), .Y(N263) );
  AO21X1TF U919 ( .A0(N325), .A1(N393), .B0(N122), .Y(N458) );
  MXI2X1TF U920 ( .A(N224), .B(N152), .S0(REG_A[15]), .Y(N260) );
  NAND2X1TF U921 ( .A(N1032), .B(N24), .Y(N231) );
  NAND2BX1TF U922 ( .AN(N238), .B(N490), .Y(N239) );
  AOI2BB1X1TF U923 ( .A0N(N1032), .A1N(N235), .B0(N182), .Y(N240) );
  OAI2BB1X1TF U924 ( .A0N(N182), .A1N(N569), .B0(N227), .Y(N228) );
  CLKBUFX2TF U925 ( .A(N1181), .Y(N222) );
  CLKBUFX2TF U926 ( .A(N1178), .Y(N221) );
  CLKBUFX2TF U927 ( .A(N378), .Y(N220) );
  OR3X1TF U928 ( .A(N542), .B(N181), .C(CODE_TYPE[3]), .Y(N540) );
  NAND2X1TF U929 ( .A(N467), .B(REG_A[12]), .Y(N746) );
  NAND2X1TF U930 ( .A(N735), .B(REG_A[10]), .Y(N744) );
  OAI221XLTF U931 ( .A0(N1130), .A1(REG_A[0]), .B0(REG_B[0]), .B1(REG_A[1]), 
        .C0(N200), .Y(N764) );
  NAND2X1TF U932 ( .A(N393), .B(REG_A[9]), .Y(N761) );
  NAND2X1TF U933 ( .A(CODE_TYPE[4]), .B(N542), .Y(N1007) );
  NAND2X1TF U934 ( .A(N467), .B(REG_A[11]), .Y(N737) );
  NAND2X1TF U935 ( .A(N467), .B(REG_A[13]), .Y(N422) );
  OAI222X1TF U936 ( .A0(N128), .A1(N386), .B0(N126), .B1(N385), .C0(N421), 
        .C1(N217), .Y(N468) );
  NAND2X1TF U937 ( .A(N735), .B(REG_A[11]), .Y(N805) );
  NAND2X1TF U938 ( .A(N777), .B(N201), .Y(N730) );
  NAND2X1TF U939 ( .A(N393), .B(REG_A[10]), .Y(N427) );
  NAND2X1TF U940 ( .A(REG_A[9]), .B(N467), .Y(N807) );
  NAND2X1TF U941 ( .A(N735), .B(REG_A[7]), .Y(N824) );
  NAND4X1TF U942 ( .A(N733), .B(N427), .C(N807), .D(N824), .Y(N872) );
  AOI222XLTF U943 ( .A0(N430), .A1(N846), .B0(N872), .B1(N848), .C0(N429), 
        .C1(N844), .Y(N432) );
  OAI222X1TF U944 ( .A0(N126), .A1(N386), .B0(N128), .B1(N384), .C0(N416), 
        .C1(N217), .Y(N4860) );
  NAND2X1TF U945 ( .A(N735), .B(REG_A[8]), .Y(N758) );
  NAND2X1TF U946 ( .A(N467), .B(REG_A[10]), .Y(N762) );
  NAND2X1TF U947 ( .A(N467), .B(REG_A[2]), .Y(N767) );
  NAND2X1TF U948 ( .A(REG_A[6]), .B(N467), .Y(N759) );
  NAND3X1TF U949 ( .A(N554), .B(START), .C(N183), .Y(N716) );
  NOR4XLTF U950 ( .A(N223), .B(N1009), .C(N875), .D(N544), .Y(N167) );
  NAND2X1TF U951 ( .A(N696), .B(I_ADDR[4]), .Y(N697) );
  NAND2X1TF U952 ( .A(N701), .B(I_ADDR[6]), .Y(N706) );
  NOR2BX1TF U953 ( .AN(N715), .B(N714), .Y(N168) );
  NAND2X1TF U954 ( .A(STATE[0]), .B(N195), .Y(N711) );
  NOR4XLTF U955 ( .A(N729), .B(N711), .C(N179), .D(N875), .Y(N616) );
  NAND2X1TF U956 ( .A(N24), .B(N569), .Y(N728) );
  NOR2BX1TF U957 ( .AN(N5170), .B(N714), .Y(N5160) );
  NAND2X1TF U958 ( .A(N546), .B(N5170), .Y(N704) );
  AO22X1TF U959 ( .A0(D_ADDR[8]), .A1(N709), .B0(I_ADDR[8]), .B1(N702), .Y(
        N536) );
  OAI221XLTF U960 ( .A0(N24), .A1(N182), .B0(N223), .B1(N391), .C0(N569), .Y(
        N539) );
  NAND2X1TF U961 ( .A(I_ADDR[1]), .B(I_ADDR[2]), .Y(N693) );
  OAI2BB2XLTF U962 ( .B0(STATE[3]), .B1(N716), .A0N(N715), .A1N(N714), .Y(N717) );
  NAND2X1TF U963 ( .A(N210), .B(N724), .Y(N1018) );
  NAND2X1TF U964 ( .A(N182), .B(N1032), .Y(N1003) );
  NAND2X1TF U965 ( .A(N864), .B(REG_B[3]), .Y(N778) );
  NAND2X1TF U966 ( .A(N393), .B(REG_A[15]), .Y(N792) );
  NAND2X1TF U967 ( .A(N864), .B(N846), .Y(N834) );
  NAND2X1TF U968 ( .A(N387), .B(N846), .Y(N869) );
  NAND4X1TF U969 ( .A(N759), .B(N758), .C(N757), .D(N756), .Y(N841) );
  AOI222XLTF U970 ( .A0(N841), .A1(N848), .B0(N837), .B1(N846), .C0(N763), 
        .C1(N844), .Y(N770) );
  AOI2BB2X1TF U971 ( .B0(REG_A[3]), .B1(N795), .A0N(N204), .A1N(N794), .Y(N796) );
  NAND4BX1TF U972 ( .AN(N813), .B(N807), .C(N806), .D(N805), .Y(N847) );
  AOI222XLTF U973 ( .A0(N849), .A1(N848), .B0(N847), .B1(N846), .C0(N845), 
        .C1(N844), .Y(N858) );
  NAND2X1TF U974 ( .A(N204), .B(N864), .Y(N866) );
  NAND2X1TF U975 ( .A(N1012), .B(N908), .Y(N1177) );
  AOI2BB2X1TF U976 ( .B0(IO_DATAINA[2]), .B1(N169), .A0N(N380), .A1N(N128), 
        .Y(N1064) );
  NAND3X1TF U977 ( .A(N1122), .B(N1121), .C(N1120), .Y(N491) );
  AO22X1TF U978 ( .A0(N1188), .A1(N199), .B0(N1189), .B1(I_DATAIN[4]), .Y(N523) );
endmodule


module SCPU_SRAM_8BIT_ALU_SPI_TOP_VG ( CLK, RST_N, CTRL_MODE, CTRL_BGN, CPU_BGN, 
        LOAD_N, CTRL_SI, ADC_PI, CTRL_RDY, CTRL_SO, NXT, SCLK1, SCLK2, LAT, 
        SPI_SO );
  input [1:0] CTRL_MODE;
  input [9:0] ADC_PI;
  output [1:0] NXT;
  input CLK, RST_N, CTRL_BGN, CPU_BGN, LOAD_N, CTRL_SI;
  output CTRL_RDY, CTRL_SO, SCLK1, SCLK2, LAT, SPI_SO;
  wire   CEN_AFTER_MUX, WEN_AFTER_MUX, I_CLK, I_RST_N, I_CTRL_BGN, I_CPU_BGN,
         I_LOAD_N, I_CTRL_SI, I_CTRL_SO, I_SCLK1, I_SCLK2, I_SPI_SO,
         SCPU_CTRL_SPI_CEN, \SCPU_CTRL_SPI_IO_DATAOUTB[0] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[1] , \SCPU_CTRL_SPI_IO_DATAOUTB[2] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[3] , \SCPU_CTRL_SPI_IO_DATAOUTB[4] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[5] , \SCPU_CTRL_SPI_IO_DATAOUTB[6] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[7] , \SCPU_CTRL_SPI_IO_DATAOUTB[8] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[9] , \SCPU_CTRL_SPI_IO_DATAOUTB[10] ,
         \SCPU_CTRL_SPI_IO_DATAOUTB[11] , \SCPU_CTRL_SPI_IO_DATAOUTB[12] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[0] , \SCPU_CTRL_SPI_IO_DATAOUTA[1] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[2] , \SCPU_CTRL_SPI_IO_DATAOUTA[3] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[4] , \SCPU_CTRL_SPI_IO_DATAOUTA[5] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[6] , \SCPU_CTRL_SPI_IO_DATAOUTA[7] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[8] , \SCPU_CTRL_SPI_IO_DATAOUTA[9] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[10] , \SCPU_CTRL_SPI_IO_DATAOUTA[11] ,
         \SCPU_CTRL_SPI_IO_DATAOUTA[12] , \SCPU_CTRL_SPI_IO_CONTROL[0] ,
         \SCPU_CTRL_SPI_IO_CONTROL[1] , \SCPU_CTRL_SPI_IO_CONTROL[2] ,
         \SCPU_CTRL_SPI_IO_CONTROL[3] , \SCPU_CTRL_SPI_IO_CONTROL[4] ,
         \SCPU_CTRL_SPI_IO_CONTROL[5] , \SCPU_CTRL_SPI_IO_CONTROL[6] ,
         SCPU_CTRL_SPI_D_WE, SCPU_CTRL_SPI_IS_I_ADDR, SCPU_CTRL_SPI_CCT_N57,
         SCPU_CTRL_SPI_CCT_N56, SCPU_CTRL_SPI_CCT_N55, SCPU_CTRL_SPI_CCT_N53,
         SCPU_CTRL_SPI_CCT_N52, SCPU_CTRL_SPI_CCT_N51,
         SCPU_CTRL_SPI_CCT_IS_SHIFT, \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[3] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[5] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ,
         \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[7] , \SCPU_CTRL_SPI_CCT_REG_BITS[1] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[2] , \SCPU_CTRL_SPI_CCT_REG_BITS[3] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[4] , \SCPU_CTRL_SPI_CCT_REG_BITS[5] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[6] , \SCPU_CTRL_SPI_CCT_REG_BITS[7] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[8] , \SCPU_CTRL_SPI_CCT_REG_BITS[9] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[10] , \SCPU_CTRL_SPI_CCT_REG_BITS[11] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[12] , \SCPU_CTRL_SPI_CCT_REG_BITS[13] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[14] , \SCPU_CTRL_SPI_CCT_REG_BITS[15] ,
         \SCPU_CTRL_SPI_CCT_REG_BITS[16] , \SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ,
         SCPU_CTRL_SPI_PUT_N108, SCPU_CTRL_SPI_PUT_N107,
         SCPU_CTRL_SPI_PUT_N106, \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ,
         \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ,
         \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ,
         \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ,
         \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] , \SCPU_CTRL_SPI_PUT_SPI_STATE[0] ,
         \SCPU_CTRL_SPI_PUT_SPI_STATE[1] , \SCPU_CTRL_SPI_PUT_CNT_STATE[0] ,
         \SCPU_CTRL_SPI_PUT_CNT_STATE[1] , \SCPU_CTRL_SPI_PUT_CNT_STATE[2] ,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N79, N80, N81, N82, N83, N84, N85, N86, N87, N91, N93, N101,
         N104, N158, N164, N165, N189, N190, N191, N192, N193, N194, N195,
         N196, N197, N198, N199, N200, N201, N202, N203, N204, N205, N206,
         N207, N208, N209, N210, N212, N213, N214, N215, N216, N218, N219,
         N220, N221, N222, N233, N234, N241, N271, N272, N273, N274, N275,
         N276, N277, N279, N280, N281, N282, N283, N284, N285, N286, N287,
         N288, N289, N290, N291, N292, N293, N294, N295, N296, N297, N298,
         N299, N300, N301, N302, N303, N304, N305, N306, N307, N308, N309,
         N310, N311, N312, N313, N314, N315, N316, N317, N318, N319, N320,
         N321, N322, N323, N324, N325, N326, N327, N328, N329, N330, N331,
         N332, N333, N334, N335, N336, N337, N338, N339, N340, N341, N342,
         N343, N344, N345, N346, N347, N348, N349, N350, N351, N352, N353,
         N354, N355, N356, N357, N358, N359, N360, N361, N362, N363, N364,
         N365, N366, N367, N368, N369, N370, N371, N372, N373, N374, N375,
         N376, N377, N378, N379, N380, N381, N382, N383, N384, N385, N386,
         N387, N388, N389, N390, N391, N392, N393, N394, N395, N396, N397,
         N398, N399, N400, N401, N402, N403, N404, N405, N406, N407, N408,
         N409, N410, N411, N412, N413, N414, N415, N416, N417, N418, N419,
         N420, N421, N422, N423, N424, N425, N426, N427, N428, N429, N430,
         N431;
  wire   [8:0] A_AFTER_MUX;
  wire   [7:0] D_AFTER_MUX;
  wire   [7:0] Q_FROM_SRAM;
  wire   [1:0] I_CTRL_MODE;
  wire   [9:0] I_ADC_PI;
  wire   [1:0] I_NXT;
  wire   [8:0] SCPU_CTRL_SPI_A_SPI;
  wire   [12:0] SCPU_CTRL_SPI_POUT;
  wire   [12:0] SCPU_CTRL_SPI_FOUT;
  wire   [9:0] SCPU_CTRL_SPI_IO_OFFSET;
  wire   [12:0] SCPU_CTRL_SPI_IO_DATAINA;
  wire   [0:0] SCPU_CTRL_SPI_IO_STATUS;
  wire   [7:0] SCPU_CTRL_SPI_D_DATAOUT;
  wire   [8:1] SCPU_CTRL_SPI_D_ADDR;
  wire   [8:0] SCPU_CTRL_SPI_I_ADDR;
  wire   [7:0] SCPU_CTRL_SPI_D_DATAIN;
  wire   [7:0] SCPU_CTRL_SPI_I_DATAIN;
  wire   [7:1] SCPU_CTRL_SPI_PUT_SRAM_REGS;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21;

  RA1SHD_IBM512X8 sram ( .Q(Q_FROM_SRAM), .A(A_AFTER_MUX), .D(D_AFTER_MUX), 
        .CLK(I_CLK), .CEN(CEN_AFTER_MUX), .WEN(WEN_AFTER_MUX) );
  PIC ipad_clk ( .IE(1'b1), .P(CLK), .Y(I_CLK) );
  PIC ipad_rst_n ( .IE(1'b1), .P(RST_N), .Y(I_RST_N) );
  PIC ipad_ctrl_mode0 ( .IE(1'b1), .P(CTRL_MODE[0]), .Y(I_CTRL_MODE[0]) );
  PIC ipad_ctrl_mode1 ( .IE(1'b1), .P(CTRL_MODE[1]), .Y(I_CTRL_MODE[1]) );
  PIC ipad_ctrl_bgn ( .IE(1'b1), .P(CTRL_BGN), .Y(I_CTRL_BGN) );
  PIC ipad_cpu_str ( .IE(1'b1), .P(CPU_BGN), .Y(I_CPU_BGN) );
  PIC ipad_load_n ( .IE(1'b1), .P(LOAD_N), .Y(I_LOAD_N) );
  PIC ipad_ctrl_si ( .IE(1'b1), .P(CTRL_SI), .Y(I_CTRL_SI) );
  PIC ipad_adc_pi0 ( .IE(1'b1), .P(ADC_PI[0]), .Y(I_ADC_PI[0]) );
  PIC ipad_adc_pi1 ( .IE(1'b1), .P(ADC_PI[1]), .Y(I_ADC_PI[1]) );
  PIC ipad_adc_pi2 ( .IE(1'b1), .P(ADC_PI[2]), .Y(I_ADC_PI[2]) );
  PIC ipad_adc_pi3 ( .IE(1'b1), .P(ADC_PI[3]), .Y(I_ADC_PI[3]) );
  PIC ipad_adc_pi4 ( .IE(1'b1), .P(ADC_PI[4]), .Y(I_ADC_PI[4]) );
  PIC ipad_adc_pi5 ( .IE(1'b1), .P(ADC_PI[5]), .Y(I_ADC_PI[5]) );
  PIC ipad_adc_pi6 ( .IE(1'b1), .P(ADC_PI[6]), .Y(I_ADC_PI[6]) );
  PIC ipad_adc_pi7 ( .IE(1'b1), .P(ADC_PI[7]), .Y(I_ADC_PI[7]) );
  PIC ipad_adc_pi8 ( .IE(1'b1), .P(ADC_PI[8]), .Y(I_ADC_PI[8]) );
  PIC ipad_adc_pi9 ( .IE(1'b1), .P(ADC_PI[9]), .Y(I_ADC_PI[9]) );
  POC8B opad_ctrl_rdy ( .A(N220), .P(CTRL_RDY) );
  POC8B opad_ctrl_so ( .A(I_CTRL_SO), .P(CTRL_SO) );
  POC8B opad_nxt0 ( .A(I_NXT[0]), .P(NXT[0]) );
  POC8B opad_nxt1 ( .A(I_NXT[1]), .P(NXT[1]) );
  POC8B opad_sclk1 ( .A(I_SCLK1), .P(SCLK1) );
  POC8B opad_sclk2 ( .A(I_SCLK2), .P(SCLK2) );
  POC8B opad_lat ( .A(N222), .P(LAT) );
  POC8B opad_spi_so ( .A(I_SPI_SO), .P(SPI_SO) );
  SHARE_SUPERALU_VG \scpu_ctrl_spi/ALU_01  ( .CLK(I_CLK), .RST_N(I_RST_N), .X_IN(
        {\SCPU_CTRL_SPI_IO_DATAOUTA[12] , \SCPU_CTRL_SPI_IO_DATAOUTA[11] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[10] , \SCPU_CTRL_SPI_IO_DATAOUTA[9] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[8] , \SCPU_CTRL_SPI_IO_DATAOUTA[7] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[6] , \SCPU_CTRL_SPI_IO_DATAOUTA[5] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[4] , \SCPU_CTRL_SPI_IO_DATAOUTA[3] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[2] , \SCPU_CTRL_SPI_IO_DATAOUTA[1] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[0] }), .Y_IN({
        \SCPU_CTRL_SPI_IO_DATAOUTB[12] , \SCPU_CTRL_SPI_IO_DATAOUTB[11] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[10] , \SCPU_CTRL_SPI_IO_DATAOUTB[9] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[8] , \SCPU_CTRL_SPI_IO_DATAOUTB[7] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[6] , \SCPU_CTRL_SPI_IO_DATAOUTB[5] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[4] , \SCPU_CTRL_SPI_IO_DATAOUTB[3] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[2] , \SCPU_CTRL_SPI_IO_DATAOUTB[1] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[0] }), .ALU_START(N272), .ALU_TYPE({
        \SCPU_CTRL_SPI_IO_CONTROL[4] , \SCPU_CTRL_SPI_IO_CONTROL[3] , 
        \SCPU_CTRL_SPI_IO_CONTROL[2] }), .MODE_TYPE({
        \SCPU_CTRL_SPI_IO_CONTROL[1] , \SCPU_CTRL_SPI_IO_CONTROL[0] }), 
        .OFFSET(SCPU_CTRL_SPI_IO_OFFSET), .FOUT(SCPU_CTRL_SPI_FOUT), .POUT(
        SCPU_CTRL_SPI_POUT), .ALU_IS_DONE(SCPU_CTRL_SPI_IO_STATUS[0]) );
  SERIAL_CPU_8BIT_VG \scpu_ctrl_spi/uut  ( .CLK(I_CLK), .ENABLE(1'b0), .RST_N(
        I_RST_N), .START(I_CPU_BGN), .I_DATAIN(SCPU_CTRL_SPI_I_DATAIN), 
        .D_DATAIN(SCPU_CTRL_SPI_D_DATAIN), .IS_I_ADDR(SCPU_CTRL_SPI_IS_I_ADDR), 
        .NXT(I_NXT), .I_ADDR(SCPU_CTRL_SPI_I_ADDR), .D_ADDR({
        SCPU_CTRL_SPI_D_ADDR, SYNOPSYS_UNCONNECTED__0}), .D_WE(
        SCPU_CTRL_SPI_D_WE), .D_DATAOUT(SCPU_CTRL_SPI_D_DATAOUT), .IO_STATUS({
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, N221, SCPU_CTRL_SPI_IO_STATUS[0]}), .IO_CONTROL({
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, \SCPU_CTRL_SPI_IO_CONTROL[6] , 
        \SCPU_CTRL_SPI_IO_CONTROL[5] , \SCPU_CTRL_SPI_IO_CONTROL[4] , 
        \SCPU_CTRL_SPI_IO_CONTROL[3] , \SCPU_CTRL_SPI_IO_CONTROL[2] , 
        \SCPU_CTRL_SPI_IO_CONTROL[1] , \SCPU_CTRL_SPI_IO_CONTROL[0] }), 
        .IO_DATAINA({1'b0, 1'b0, 1'b0, SCPU_CTRL_SPI_IO_DATAINA}), 
        .IO_DATAINB({1'b0, 1'b0, 1'b0, SCPU_CTRL_SPI_POUT}), .IO_DATAOUTA({
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, \SCPU_CTRL_SPI_IO_DATAOUTA[12] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[11] , \SCPU_CTRL_SPI_IO_DATAOUTA[10] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[9] , \SCPU_CTRL_SPI_IO_DATAOUTA[8] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[7] , \SCPU_CTRL_SPI_IO_DATAOUTA[6] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[5] , \SCPU_CTRL_SPI_IO_DATAOUTA[4] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[3] , \SCPU_CTRL_SPI_IO_DATAOUTA[2] , 
        \SCPU_CTRL_SPI_IO_DATAOUTA[1] , \SCPU_CTRL_SPI_IO_DATAOUTA[0] }), 
        .IO_DATAOUTB({SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, \SCPU_CTRL_SPI_IO_DATAOUTB[12] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[11] , \SCPU_CTRL_SPI_IO_DATAOUTB[10] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[9] , \SCPU_CTRL_SPI_IO_DATAOUTB[8] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[7] , \SCPU_CTRL_SPI_IO_DATAOUTB[6] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[5] , \SCPU_CTRL_SPI_IO_DATAOUTB[4] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[3] , \SCPU_CTRL_SPI_IO_DATAOUTB[2] , 
        \SCPU_CTRL_SPI_IO_DATAOUTB[1] , \SCPU_CTRL_SPI_IO_DATAOUTB[0] }), 
        .IO_OFFSET({SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SCPU_CTRL_SPI_IO_OFFSET}) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[7]  ( .D(N158), .RN(
        SCPU_CTRL_SPI_CCT_N57), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[7] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[5]  ( .D(N158), .RN(
        SCPU_CTRL_SPI_CCT_N55), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[5] ), .QN(N292) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[3]  ( .D(N158), .RN(
        SCPU_CTRL_SPI_CCT_N53), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[3] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[2]  ( .D(N158), .RN(
        SCPU_CTRL_SPI_CCT_N52), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[1]  ( .D(N158), .RN(
        SCPU_CTRL_SPI_CCT_N51), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ) );
  DFFTRX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[6]  ( .D(N158), .RN(
        SCPU_CTRL_SPI_CCT_N56), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ) );
  DFFRX2TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[3]  ( .D(N208), .CK(I_CLK), 
        .RN(N273), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ), .QN(N294) );
  DFFRX2TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[0]  ( .D(N205), .CK(I_CLK), 
        .RN(N274), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .QN(N291) );
  DFFRX2TF \scpu_ctrl_spi/put/spi_state_reg[2]  ( .D(N212), .CK(I_CLK), .RN(
        N274), .Q(N289), .QN(N101) );
  DFFRX2TF \scpu_ctrl_spi/put/cnt_state_reg[1]  ( .D(SCPU_CTRL_SPI_PUT_N107), 
        .CK(I_CLK), .RN(N274), .Q(\SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .QN(N288)
         );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[4]  ( .D(N45), .CK(I_CLK), 
        .SN(N44), .RN(N43), .QN(N285) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[0]  ( .D(N33), .CK(I_CLK), 
        .SN(N32), .RN(N31), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .QN(N284)
         );
  DFFRX2TF \scpu_ctrl_spi/put/spi_state_reg[1]  ( .D(N210), .CK(I_CLK), .RN(
        N274), .Q(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .QN(N283) );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[3]  ( .D(N42), .CK(I_CLK), 
        .SN(N41), .RN(N40), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] ), .QN(N282)
         );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[2]  ( .D(N39), .CK(I_CLK), 
        .SN(N38), .RN(N37), .QN(N281) );
  DFFSX2TF \scpu_ctrl_spi/put/cnt_state_reg[0]  ( .D(SCPU_CTRL_SPI_PUT_N106), 
        .CK(I_CLK), .SN(N274), .Q(\SCPU_CTRL_SPI_PUT_CNT_STATE[0] ), .QN(N280)
         );
  DFFSRX2TF \scpu_ctrl_spi/put/cnt_addr_len_reg[1]  ( .D(N36), .CK(I_CLK), 
        .SN(N35), .RN(N34), .Q(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ), .QN(N279)
         );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[7]  ( .D(N189), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[7] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[6]  ( .D(N190), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[6] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[5]  ( .D(N191), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[5] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[4]  ( .D(N192), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[4] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[3]  ( .D(N193), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[3] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[2]  ( .D(N194), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[2] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[1]  ( .D(N195), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[1] ) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[7]  ( .D(N204), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[7]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[6]  ( .D(N198), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[6]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[5]  ( .D(N199), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[5]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[4]  ( .D(N200), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[4]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[3]  ( .D(N201), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[3]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[2]  ( .D(N202), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[2]) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[1]  ( .D(N203), .CK(I_CLK), .Q(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[1]) );
  DFFTRX1TF \scpu_ctrl_spi/cct/is_shift_reg  ( .D(N164), .RN(N165), .CK(I_CLK), 
        .QN(SCPU_CTRL_SPI_CCT_IS_SHIFT) );
  DFFQX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[4]  ( .D(N215), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/cnt_bit_load_reg[0]  ( .D(N214), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ) );
  DFFQX1TF \scpu_ctrl_spi/put/sram_regs_reg[0]  ( .D(N197), .CK(I_CLK), .Q(
        I_SPI_SO) );
  DFFQX1TF \scpu_ctrl_spi/cct/reg_bits_reg[0]  ( .D(N196), .CK(I_CLK), .Q(
        I_CTRL_SO) );
  DFFNSRX4TF \scpu_ctrl_spi/put/spi_MUX_reg  ( .D(N213), .CKN(I_CLK), .SN(1'b1), .RN(1'b1), .Q(N305), .QN(N104) );
  DFFNSRXLTF \scpu_ctrl_spi/cct/D_WE_reg  ( .D(N218), .CKN(I_CLK), .SN(1'b1), 
        .RN(1'b1), .QN(N287) );
  DFFNSRX1TF \scpu_ctrl_spi/put/sram_addr_reg[7]  ( .D(N86), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[7]), .QN(N290) );
  DFFNSRXLTF \scpu_ctrl_spi/cct/CEN_reg  ( .D(N219), .CKN(I_CLK), .SN(1'b1), 
        .RN(1'b1), .Q(SCPU_CTRL_SPI_CEN) );
  DFFNSRXLTF \scpu_ctrl_spi/put/sram_addr_reg[8]  ( .D(N87), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[8]) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[15]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[16] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[15] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[14]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[15] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[14] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[13]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[14] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[13] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[12]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[13] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[12] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[11]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[12] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[11] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[10]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[11] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[10] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[9]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[10] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[9] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[8]  ( .D(
        \SCPU_CTRL_SPI_CCT_REG_BITS[9] ), .E(N241), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_REG_BITS[8] ) );
  EDFFX1TF \scpu_ctrl_spi/cct/reg_bits_reg[16]  ( .D(I_CTRL_SI), .E(N241), 
        .CK(I_CLK), .Q(\SCPU_CTRL_SPI_CCT_REG_BITS[16] ) );
  DFFQX1TF \scpu_ctrl_spi/cct/ctrl_state_reg[0]  ( .D(N216), .CK(I_CLK), .Q(
        \SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ) );
  EDFFTRXLTF \scpu_ctrl_spi/cct/ctrl_state_reg[1]  ( .RN(I_CTRL_BGN), .D(1'b1), 
        .E(N234), .CK(I_CLK), .Q(N286), .QN(N93) );
  DFFRX1TF \scpu_ctrl_spi/put/spi_state_reg[0]  ( .D(N209), .CK(I_CLK), .RN(
        \SCPU_CTRL_SPI_IO_CONTROL[6] ), .Q(\SCPU_CTRL_SPI_PUT_SPI_STATE[0] )
         );
  DFFRX1TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[1]  ( .D(N206), .CK(I_CLK), 
        .RN(N274), .Q(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ) );
  DFFRX1TF \scpu_ctrl_spi/put/cnt_state_reg[2]  ( .D(SCPU_CTRL_SPI_PUT_N108), 
        .CK(I_CLK), .RN(N274), .Q(\SCPU_CTRL_SPI_PUT_CNT_STATE[2] ) );
  DFFRX1TF \scpu_ctrl_spi/put/cnt_bit_sent_reg[2]  ( .D(N207), .CK(I_CLK), 
        .RN(\SCPU_CTRL_SPI_IO_CONTROL[6] ), .Q(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[1]  ( .D(N80), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[1]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[3]  ( .D(N82), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[3]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[5]  ( .D(N84), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[5]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[2]  ( .D(N81), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[2]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[6]  ( .D(N85), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[6]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[4]  ( .D(N83), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[4]) );
  DFFNSRX2TF \scpu_ctrl_spi/put/sram_addr_reg[0]  ( .D(N79), .CKN(I_CLK), .SN(
        1'b1), .RN(1'b1), .Q(SCPU_CTRL_SPI_A_SPI[0]), .QN(N293) );
  NOR2BX1TF U243 ( .AN(SCPU_CTRL_SPI_FOUT[10]), .B(N271), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[10]) );
  NOR2BX1TF U244 ( .AN(SCPU_CTRL_SPI_FOUT[11]), .B(N271), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[11]) );
  NOR2BX1TF U245 ( .AN(SCPU_CTRL_SPI_FOUT[12]), .B(N295), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[12]) );
  AO21X1TF U246 ( .A0(N279), .A1(N427), .B0(N281), .Y(N233) );
  OAI21X1TF U247 ( .A0(N429), .A1(N430), .B0(N233), .Y(N39) );
  OA21XLTF U248 ( .A0(N275), .A1(I_CTRL_MODE[0]), .B0(N328), .Y(N234) );
  CLKBUFX2TF U249 ( .A(N91), .Y(N241) );
  INVX2TF U263 ( .A(N295), .Y(N272) );
  CLKBUFX2TF U264 ( .A(\SCPU_CTRL_SPI_CCT_CTRL_STATE[0] ), .Y(N275) );
  NAND2XLTF U265 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[0] ), .B(N296), .Y(N32) );
  NAND2XLTF U266 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[1] ), .B(N296), .Y(N35) );
  NAND2XLTF U267 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[4] ), .B(N296), .Y(N44) );
  NAND2XLTF U268 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[2] ), .B(N296), .Y(N38) );
  NAND2XLTF U269 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[3] ), .B(N296), .Y(N41) );
  INVX1TF U270 ( .A(N408), .Y(N411) );
  NOR3BX1TF U271 ( .AN(SCPU_CTRL_SPI_CCT_IS_SHIFT), .B(N286), .C(N373), .Y(N91) );
  INVX2TF U272 ( .A(N296), .Y(N273) );
  INVX2TF U273 ( .A(N275), .Y(N373) );
  NOR3X1TF U274 ( .A(N275), .B(N286), .C(N327), .Y(N330) );
  NAND2XLTF U275 ( .A(N340), .B(N395), .Y(N339) );
  INVX2TF U276 ( .A(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .Y(N295) );
  NOR2X4TF U277 ( .A(SCPU_CTRL_SPI_CEN), .B(N327), .Y(N325) );
  NAND2XLTF U278 ( .A(SCPU_CTRL_SPI_A_SPI[0]), .B(SCPU_CTRL_SPI_A_SPI[1]), .Y(
        N421) );
  OR2X2TF U279 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ), .B(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .Y(N300) );
  INVX2TF U280 ( .A(\SCPU_CTRL_SPI_IO_CONTROL[6] ), .Y(N296) );
  INVX2TF U281 ( .A(N272), .Y(N271) );
  INVX2TF U282 ( .A(N296), .Y(N274) );
  NOR3X4TF U283 ( .A(I_CTRL_BGN), .B(N298), .C(N361), .Y(N370) );
  NAND4BX2TF U284 ( .AN(N219), .B(I_CTRL_BGN), .C(SCPU_CTRL_SPI_CCT_IS_SHIFT), 
        .D(N374), .Y(N384) );
  INVX2TF U285 ( .A(I_CTRL_BGN), .Y(N276) );
  CLKBUFX2TF U286 ( .A(N241), .Y(N297) );
  NOR3X4TF U287 ( .A(N360), .B(N359), .C(N298), .Y(N371) );
  NOR3X2TF U288 ( .A(\SCPU_CTRL_SPI_PUT_CNT_STATE[0] ), .B(
        \SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .C(\SCPU_CTRL_SPI_PUT_CNT_STATE[2] ), .Y(N395) );
  INVX2TF U289 ( .A(N429), .Y(N277) );
  NOR2BX1TF U290 ( .AN(N344), .B(N428), .Y(N426) );
  INVX2TF U291 ( .A(I_CTRL_BGN), .Y(N327) );
  NOR2X1TF U292 ( .A(N348), .B(N362), .Y(N358) );
  NAND2X1TF U293 ( .A(I_CTRL_BGN), .B(N329), .Y(N337) );
  NOR2X1TF U294 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[3] ), .B(N301), .Y(N164)
         );
  AOI222XLTF U295 ( .A0(N371), .A1(I_SPI_SO), .B0(N370), .B1(Q_FROM_SRAM[0]), 
        .C0(SCPU_CTRL_SPI_PUT_SRAM_REGS[1]), .C1(N369), .Y(N372) );
  AOI222XLTF U296 ( .A0(N371), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[3]), .B0(N370), 
        .B1(Q_FROM_SRAM[3]), .C0(N369), .C1(SCPU_CTRL_SPI_PUT_SRAM_REGS[4]), 
        .Y(N365) );
  AOI222XLTF U297 ( .A0(N371), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[2]), .B0(N370), 
        .B1(Q_FROM_SRAM[2]), .C0(N369), .C1(SCPU_CTRL_SPI_PUT_SRAM_REGS[3]), 
        .Y(N364) );
  AOI222XLTF U298 ( .A0(N371), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[1]), .B0(N370), 
        .B1(Q_FROM_SRAM[1]), .C0(N369), .C1(SCPU_CTRL_SPI_PUT_SRAM_REGS[2]), 
        .Y(N363) );
  AOI222XLTF U299 ( .A0(N371), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[5]), .B0(N370), 
        .B1(Q_FROM_SRAM[5]), .C0(N369), .C1(SCPU_CTRL_SPI_PUT_SRAM_REGS[6]), 
        .Y(N367) );
  AOI222XLTF U300 ( .A0(N371), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[4]), .B0(N370), 
        .B1(Q_FROM_SRAM[4]), .C0(N369), .C1(SCPU_CTRL_SPI_PUT_SRAM_REGS[5]), 
        .Y(N366) );
  AOI222XLTF U301 ( .A0(N371), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[6]), .B0(
        SCPU_CTRL_SPI_PUT_SRAM_REGS[7]), .B1(N369), .C0(N370), .C1(
        Q_FROM_SRAM[6]), .Y(N368) );
  NOR2X1TF U302 ( .A(N346), .B(N101), .Y(N359) );
  NAND2X1TF U303 ( .A(N319), .B(N318), .Y(A_AFTER_MUX[7]) );
  NAND2X1TF U304 ( .A(N315), .B(N314), .Y(A_AFTER_MUX[5]) );
  NAND2X1TF U305 ( .A(N311), .B(N310), .Y(A_AFTER_MUX[3]) );
  NAND2X1TF U306 ( .A(N309), .B(N308), .Y(A_AFTER_MUX[2]) );
  CLKBUFX2TF U307 ( .A(N296), .Y(N298) );
  NAND2X1TF U308 ( .A(N338), .B(N101), .Y(N428) );
  NOR2X1TF U309 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ), .B(N302), .Y(N303)
         );
  NAND2X1TF U310 ( .A(N292), .B(N332), .Y(N302) );
  NOR2X1TF U311 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ), .B(N333), .Y(N332)
         );
  OAI2BB2XLTF U312 ( .B0(N398), .B1(N397), .A0N(
        \SCPU_CTRL_SPI_PUT_CNT_STATE[2] ), .A1N(N396), .Y(
        SCPU_CTRL_SPI_PUT_N108) );
  NOR2X1TF U313 ( .A(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ), .B(N343), .Y(N348)
         );
  NAND2X1TF U314 ( .A(N164), .B(N165), .Y(N329) );
  OR3X1TF U315 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ), .B(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ), .C(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .Y(N301) );
  NOR2X2TF U316 ( .A(N298), .B(N362), .Y(N369) );
  NOR2X1TF U317 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .B(N283), .Y(N340) );
  NAND3X1TF U318 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .B(
        \SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .C(N101), .Y(N361) );
  NOR2BX1TF U319 ( .AN(N347), .B(N101), .Y(N222) );
  AND2X2TF U320 ( .A(N325), .B(N287), .Y(N326) );
  OAI2BB1X1TF U321 ( .A0N(N325), .A1N(\SCPU_CTRL_SPI_CCT_REG_BITS[8] ), .B0(
        N304), .Y(A_AFTER_MUX[0]) );
  NAND2X1TF U322 ( .A(N324), .B(N323), .Y(A_AFTER_MUX[8]) );
  NAND2X1TF U323 ( .A(N317), .B(N316), .Y(A_AFTER_MUX[6]) );
  NAND2X1TF U324 ( .A(N313), .B(N312), .Y(A_AFTER_MUX[4]) );
  NAND2X1TF U325 ( .A(N307), .B(N306), .Y(A_AFTER_MUX[1]) );
  NOR2X2TF U326 ( .A(N385), .B(N305), .Y(N322) );
  OR2X2TF U327 ( .A(SCPU_CTRL_SPI_IS_I_ADDR), .B(I_CTRL_BGN), .Y(N385) );
  NOR2X2TF U328 ( .A(N305), .B(N393), .Y(N320) );
  NAND2X2TF U329 ( .A(SCPU_CTRL_SPI_IS_I_ADDR), .B(N327), .Y(N393) );
  NOR2X2TF U330 ( .A(I_CTRL_BGN), .B(N104), .Y(N321) );
  NAND2X1TF U331 ( .A(N275), .B(N286), .Y(N219) );
  AO22X1TF U332 ( .A0(N272), .A1(SCPU_CTRL_SPI_FOUT[8]), .B0(N295), .B1(
        I_ADC_PI[8]), .Y(SCPU_CTRL_SPI_IO_DATAINA[8]) );
  AO22X1TF U333 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[4]), .B0(N295), .B1(I_ADC_PI[4]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[4]) );
  AO22X1TF U334 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[9]), .B0(N271), .B1(I_ADC_PI[9]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[9]) );
  NAND2X1TF U335 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .B(N283), .Y(N342) );
  AO22X1TF U336 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[7]), .B0(N295), .B1(I_ADC_PI[7]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[7]) );
  AO22X1TF U337 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[6]), .B0(N295), .B1(I_ADC_PI[6]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[6]) );
  OR2X2TF U338 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[3] ), .B(
        \SCPU_CTRL_SPI_IO_CONTROL[6] ), .Y(N40) );
  OR2X2TF U339 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[0] ), .B(
        \SCPU_CTRL_SPI_IO_CONTROL[6] ), .Y(N31) );
  OR2X2TF U340 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[1] ), .B(N274), .Y(N34) );
  OR2X2TF U341 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[2] ), .B(
        \SCPU_CTRL_SPI_IO_CONTROL[6] ), .Y(N37) );
  OR2X2TF U342 ( .A(\SCPU_CTRL_SPI_IO_DATAOUTB[4] ), .B(N274), .Y(N43) );
  NOR2X1TF U343 ( .A(\SCPU_CTRL_SPI_PUT_CNT_STATE[0] ), .B(N395), .Y(
        SCPU_CTRL_SPI_PUT_N106) );
  AOI21X1TF U344 ( .A0(N431), .A1(N282), .B0(N285), .Y(N45) );
  OAI31X1TF U345 ( .A0(N351), .A1(N342), .A2(N344), .B0(N341), .Y(N212) );
  AOI32X1TF U346 ( .A0(N395), .A1(N101), .A2(N340), .B0(N289), .B1(N339), .Y(
        N341) );
  OAI21X1TF U347 ( .A0(N351), .A1(N350), .B0(N349), .Y(N209) );
  OAI21X1TF U348 ( .A0(N289), .A1(N397), .B0(\SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), 
        .Y(N349) );
  AOI211X1TF U349 ( .A0(N348), .A1(N289), .B0(N347), .C0(N277), .Y(N350) );
  OAI21X1TF U350 ( .A0(N332), .A1(N292), .B0(N302), .Y(SCPU_CTRL_SPI_CCT_N55)
         );
  AOI22X1TF U351 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .A1(N277), .B0(
        N429), .B1(N284), .Y(N33) );
  OAI32X1TF U352 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[3] ), .A1(N430), .A2(
        N429), .B0(N431), .B1(N282), .Y(N42) );
  NOR2X1TF U353 ( .A(N428), .B(N430), .Y(N431) );
  OAI32X1TF U354 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[1] ), .A1(
        \SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .A2(N429), .B0(N427), .B1(N279), 
        .Y(N36) );
  NOR2X1TF U355 ( .A(N101), .B(N351), .Y(N345) );
  AOI21X1TF U356 ( .A0(N289), .A1(N346), .B0(N395), .Y(N351) );
  NOR2X1TF U357 ( .A(\SCPU_CTRL_SPI_PUT_CNT_ADDR_LEN[0] ), .B(N428), .Y(N427)
         );
  OAI211X1TF U358 ( .A0(N358), .A1(N291), .B0(N361), .C0(N357), .Y(N205) );
  INVX2TF U359 ( .A(N337), .Y(N158) );
  AOI22X1TF U360 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[3] ), .A1(N353), .B0(
        N354), .B1(N294), .Y(N208) );
  AOI21X1TF U361 ( .A0(N359), .A1(N343), .B0(N398), .Y(N353) );
  OAI211X1TF U362 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .A1(N357), .B0(
        N361), .C0(N356), .Y(N206) );
  OAI21X1TF U363 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .A1(N398), .B0(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .Y(N356) );
  OAI22X1TF U364 ( .A0(I_CTRL_MODE[0]), .A1(N335), .B0(N334), .B1(N337), .Y(
        N215) );
  AOI21X1TF U365 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ), .A1(N333), .B0(
        N332), .Y(N334) );
  INVX2TF U366 ( .A(N164), .Y(N333) );
  INVX2TF U367 ( .A(N395), .Y(N397) );
  OAI31X1TF U368 ( .A0(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .A1(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .A2(N398), .B0(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ), .Y(N355) );
  NOR2X1TF U369 ( .A(N360), .B(N358), .Y(N398) );
  INVX2TF U370 ( .A(N352), .Y(N343) );
  NOR3X1TF U371 ( .A(\SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[2] ), .B(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[1] ), .C(
        \SCPU_CTRL_SPI_PUT_CNT_BIT_SENT[0] ), .Y(N352) );
  OAI21X1TF U372 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .A1(N337), .B0(
        N336), .Y(N214) );
  INVX2TF U373 ( .A(N331), .Y(N335) );
  NOR3BX1TF U374 ( .AN(N330), .B(I_LOAD_N), .C(N329), .Y(N331) );
  NOR4X1TF U375 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[7] ), .B(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ), .C(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[5] ), .D(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[4] ), .Y(N165) );
  INVX2TF U376 ( .A(N372), .Y(N197) );
  INVX2TF U377 ( .A(N365), .Y(N201) );
  INVX2TF U378 ( .A(N364), .Y(N202) );
  INVX2TF U379 ( .A(N363), .Y(N203) );
  INVX2TF U380 ( .A(N367), .Y(N199) );
  INVX2TF U381 ( .A(N366), .Y(N200) );
  INVX2TF U382 ( .A(N368), .Y(N198) );
  INVX2TF U383 ( .A(N359), .Y(N362) );
  INVX2TF U384 ( .A(N340), .Y(N346) );
  INVX2TF U385 ( .A(N361), .Y(N360) );
  OAI21X1TF U386 ( .A0(N389), .A1(N384), .B0(N378), .Y(N193) );
  AOI22X1TF U387 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[4] ), .A1(N297), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[3] ), .B1(N382), .Y(N378) );
  OAI21X1TF U388 ( .A0(N388), .A1(N384), .B0(N377), .Y(N194) );
  AOI22X1TF U389 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[3] ), .A1(N297), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[2] ), .B1(N382), .Y(N377) );
  OAI21X1TF U390 ( .A0(N387), .A1(N384), .B0(N376), .Y(N195) );
  AOI22X1TF U391 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[2] ), .A1(N297), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[1] ), .B1(N382), .Y(N376) );
  OAI21X1TF U392 ( .A0(N394), .A1(N384), .B0(N383), .Y(N189) );
  AOI22X1TF U393 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[8] ), .A1(N297), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[7] ), .B1(N382), .Y(N383) );
  OAI21X1TF U394 ( .A0(N391), .A1(N384), .B0(N380), .Y(N191) );
  AOI22X1TF U395 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[6] ), .A1(N297), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[5] ), .B1(N382), .Y(N380) );
  OAI21X1TF U396 ( .A0(N392), .A1(N384), .B0(N381), .Y(N190) );
  AOI22X1TF U397 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[7] ), .A1(N297), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[6] ), .B1(N382), .Y(N381) );
  OAI21X1TF U398 ( .A0(N390), .A1(N384), .B0(N379), .Y(N192) );
  AOI22X1TF U399 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[5] ), .A1(N297), .B0(
        \SCPU_CTRL_SPI_CCT_REG_BITS[4] ), .B1(N382), .Y(N379) );
  OAI21X1TF U400 ( .A0(N386), .A1(N384), .B0(N375), .Y(N196) );
  AOI22X1TF U401 ( .A0(\SCPU_CTRL_SPI_CCT_REG_BITS[1] ), .A1(N297), .B0(
        I_CTRL_SO), .B1(N382), .Y(N375) );
  OAI211X4TF U402 ( .A0(N93), .A1(N374), .B0(N275), .C0(
        SCPU_CTRL_SPI_CCT_IS_SHIFT), .Y(N382) );
  NOR2X1TF U403 ( .A(\SCPU_CTRL_SPI_PUT_SPI_STATE[1] ), .B(
        \SCPU_CTRL_SPI_PUT_SPI_STATE[0] ), .Y(N347) );
  NOR2X1TF U404 ( .A(N93), .B(N275), .Y(N220) );
  AOI32X1TF U405 ( .A0(N104), .A1(N327), .A2(SCPU_CTRL_SPI_D_WE), .B0(
        I_CTRL_BGN), .B1(N287), .Y(WEN_AFTER_MUX) );
  NOR2X1TF U406 ( .A(N390), .B(N393), .Y(SCPU_CTRL_SPI_I_DATAIN[4]) );
  NOR2X1TF U407 ( .A(N391), .B(N393), .Y(SCPU_CTRL_SPI_I_DATAIN[5]) );
  NOR2X1TF U408 ( .A(N387), .B(N393), .Y(SCPU_CTRL_SPI_I_DATAIN[1]) );
  NOR2X1TF U409 ( .A(N386), .B(N393), .Y(SCPU_CTRL_SPI_I_DATAIN[0]) );
  NOR2X1TF U410 ( .A(N388), .B(N393), .Y(SCPU_CTRL_SPI_I_DATAIN[2]) );
  NOR2X1TF U411 ( .A(N392), .B(N393), .Y(SCPU_CTRL_SPI_I_DATAIN[6]) );
  NOR2X1TF U412 ( .A(N394), .B(N393), .Y(SCPU_CTRL_SPI_I_DATAIN[7]) );
  NOR2X1TF U413 ( .A(N389), .B(N393), .Y(SCPU_CTRL_SPI_I_DATAIN[3]) );
  OAI32X1TF U414 ( .A0(N298), .A1(N338), .A2(N104), .B0(N428), .B1(N298), .Y(
        N213) );
  NOR2X1TF U415 ( .A(N386), .B(N385), .Y(SCPU_CTRL_SPI_D_DATAIN[0]) );
  INVX2TF U416 ( .A(Q_FROM_SRAM[0]), .Y(N386) );
  NOR2X1TF U417 ( .A(N391), .B(N385), .Y(SCPU_CTRL_SPI_D_DATAIN[5]) );
  INVX2TF U418 ( .A(Q_FROM_SRAM[5]), .Y(N391) );
  NOR2X1TF U419 ( .A(N390), .B(N385), .Y(SCPU_CTRL_SPI_D_DATAIN[4]) );
  INVX2TF U420 ( .A(Q_FROM_SRAM[4]), .Y(N390) );
  NOR2X1TF U421 ( .A(N389), .B(N385), .Y(SCPU_CTRL_SPI_D_DATAIN[3]) );
  INVX2TF U422 ( .A(Q_FROM_SRAM[3]), .Y(N389) );
  NOR2X1TF U423 ( .A(N392), .B(N385), .Y(SCPU_CTRL_SPI_D_DATAIN[6]) );
  INVX2TF U424 ( .A(Q_FROM_SRAM[6]), .Y(N392) );
  NOR2X1TF U425 ( .A(N394), .B(N385), .Y(SCPU_CTRL_SPI_D_DATAIN[7]) );
  INVX2TF U426 ( .A(Q_FROM_SRAM[7]), .Y(N394) );
  NOR2X1TF U427 ( .A(N387), .B(N385), .Y(SCPU_CTRL_SPI_D_DATAIN[1]) );
  INVX2TF U428 ( .A(Q_FROM_SRAM[1]), .Y(N387) );
  NOR2X1TF U429 ( .A(N388), .B(N385), .Y(SCPU_CTRL_SPI_D_DATAIN[2]) );
  INVX2TF U430 ( .A(Q_FROM_SRAM[2]), .Y(N388) );
  OAI31X1TF U431 ( .A0(SCPU_CTRL_SPI_A_SPI[3]), .A1(N425), .A2(N418), .B0(N417), .Y(N82) );
  AOI22X1TF U432 ( .A0(SCPU_CTRL_SPI_A_SPI[3]), .A1(N416), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[3] ), .B1(N299), .Y(N417) );
  AOI21X1TF U433 ( .A0(N277), .A1(N415), .B0(N299), .Y(N416) );
  OAI31X1TF U434 ( .A0(SCPU_CTRL_SPI_A_SPI[1]), .A1(N425), .A2(N293), .B0(N423), .Y(N80) );
  AOI22X1TF U435 ( .A0(SCPU_CTRL_SPI_A_SPI[1]), .A1(N422), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[1] ), .B1(N299), .Y(N423) );
  AOI21X1TF U436 ( .A0(N277), .A1(SCPU_CTRL_SPI_A_SPI[0]), .B0(N299), .Y(N422)
         );
  OAI31X1TF U437 ( .A0(SCPU_CTRL_SPI_A_SPI[2]), .A1(N425), .A2(N421), .B0(N420), .Y(N81) );
  AOI22X1TF U438 ( .A0(SCPU_CTRL_SPI_A_SPI[2]), .A1(N419), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[2] ), .B1(N299), .Y(N420) );
  AOI31X1TF U439 ( .A0(N277), .A1(SCPU_CTRL_SPI_A_SPI[0]), .A2(
        SCPU_CTRL_SPI_A_SPI[1]), .B0(N299), .Y(N419) );
  OAI31X1TF U440 ( .A0(SCPU_CTRL_SPI_A_SPI[4]), .A1(N425), .A2(N414), .B0(N413), .Y(N83) );
  AOI22X1TF U441 ( .A0(SCPU_CTRL_SPI_A_SPI[4]), .A1(N412), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[4] ), .B1(N299), .Y(N413) );
  AOI31X1TF U442 ( .A0(N277), .A1(N415), .A2(SCPU_CTRL_SPI_A_SPI[3]), .B0(N299), .Y(N412) );
  OAI31X1TF U443 ( .A0(SCPU_CTRL_SPI_A_SPI[6]), .A1(N425), .A2(N407), .B0(N406), .Y(N85) );
  AOI22X1TF U444 ( .A0(SCPU_CTRL_SPI_A_SPI[6]), .A1(N405), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[6] ), .B1(N298), .Y(N406) );
  AOI31X1TF U445 ( .A0(N426), .A1(N408), .A2(SCPU_CTRL_SPI_A_SPI[5]), .B0(N299), .Y(N405) );
  OAI31X1TF U446 ( .A0(SCPU_CTRL_SPI_A_SPI[5]), .A1(N425), .A2(N411), .B0(N410), .Y(N84) );
  AOI22X1TF U447 ( .A0(SCPU_CTRL_SPI_A_SPI[5]), .A1(N409), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[5] ), .B1(N298), .Y(N410) );
  AOI21X1TF U448 ( .A0(N277), .A1(N408), .B0(N299), .Y(N409) );
  AOI22X1TF U449 ( .A0(N322), .A1(SCPU_CTRL_SPI_D_ADDR[8]), .B0(N325), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[16] ), .Y(N323) );
  AOI22X1TF U450 ( .A0(SCPU_CTRL_SPI_A_SPI[8]), .A1(N321), .B0(N320), .B1(
        SCPU_CTRL_SPI_I_ADDR[8]), .Y(N324) );
  AOI22X1TF U451 ( .A0(N322), .A1(SCPU_CTRL_SPI_D_ADDR[7]), .B0(N325), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[15] ), .Y(N318) );
  AOI22X1TF U452 ( .A0(SCPU_CTRL_SPI_A_SPI[7]), .A1(N321), .B0(N320), .B1(
        SCPU_CTRL_SPI_I_ADDR[7]), .Y(N319) );
  AOI22X1TF U453 ( .A0(N322), .A1(SCPU_CTRL_SPI_D_ADDR[6]), .B0(N325), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[14] ), .Y(N316) );
  AOI22X1TF U454 ( .A0(SCPU_CTRL_SPI_A_SPI[6]), .A1(N321), .B0(N320), .B1(
        SCPU_CTRL_SPI_I_ADDR[6]), .Y(N317) );
  AOI22X1TF U455 ( .A0(N322), .A1(SCPU_CTRL_SPI_D_ADDR[5]), .B0(N325), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[13] ), .Y(N314) );
  AOI22X1TF U456 ( .A0(SCPU_CTRL_SPI_A_SPI[5]), .A1(N321), .B0(N320), .B1(
        SCPU_CTRL_SPI_I_ADDR[5]), .Y(N315) );
  AOI22X1TF U457 ( .A0(N322), .A1(SCPU_CTRL_SPI_D_ADDR[4]), .B0(N325), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[12] ), .Y(N312) );
  AOI22X1TF U458 ( .A0(SCPU_CTRL_SPI_A_SPI[4]), .A1(N321), .B0(N320), .B1(
        SCPU_CTRL_SPI_I_ADDR[4]), .Y(N313) );
  AOI22X1TF U459 ( .A0(N322), .A1(SCPU_CTRL_SPI_D_ADDR[3]), .B0(N325), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[11] ), .Y(N310) );
  AOI22X1TF U460 ( .A0(SCPU_CTRL_SPI_A_SPI[3]), .A1(N321), .B0(N320), .B1(
        SCPU_CTRL_SPI_I_ADDR[3]), .Y(N311) );
  AOI22X1TF U461 ( .A0(N322), .A1(SCPU_CTRL_SPI_D_ADDR[2]), .B0(N325), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[10] ), .Y(N308) );
  AOI22X1TF U462 ( .A0(SCPU_CTRL_SPI_A_SPI[2]), .A1(N321), .B0(N320), .B1(
        SCPU_CTRL_SPI_I_ADDR[2]), .Y(N309) );
  AOI22X1TF U463 ( .A0(N322), .A1(SCPU_CTRL_SPI_D_ADDR[1]), .B0(N325), .B1(
        \SCPU_CTRL_SPI_CCT_REG_BITS[9] ), .Y(N306) );
  AOI22X1TF U464 ( .A0(SCPU_CTRL_SPI_A_SPI[1]), .A1(N321), .B0(N320), .B1(
        SCPU_CTRL_SPI_I_ADDR[1]), .Y(N307) );
  OAI31X1TF U465 ( .A0(SCPU_CTRL_SPI_A_SPI[8]), .A1(N290), .A2(N402), .B0(N401), .Y(N87) );
  AOI22X1TF U466 ( .A0(SCPU_CTRL_SPI_A_SPI[8]), .A1(N400), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[8] ), .B1(N298), .Y(N401) );
  OAI21X1TF U467 ( .A0(SCPU_CTRL_SPI_A_SPI[7]), .A1(N425), .B0(N404), .Y(N400)
         );
  OAI21X1TF U468 ( .A0(N404), .A1(N290), .B0(N403), .Y(N86) );
  INVX2TF U469 ( .A(N418), .Y(N415) );
  OR2X2TF U470 ( .A(N219), .B(N374), .Y(N218) );
  OAI21X1TF U471 ( .A0(SCPU_CTRL_SPI_A_SPI[0]), .A1(N425), .B0(N424), .Y(N79)
         );
  AOI32X1TF U472 ( .A0(SCPU_CTRL_SPI_A_SPI[0]), .A1(N274), .A2(N429), .B0(
        \SCPU_CTRL_SPI_IO_DATAOUTA[0] ), .B1(N298), .Y(N424) );
  INVX2TF U473 ( .A(N426), .Y(N429) );
  NAND2X2TF U474 ( .A(N426), .B(N273), .Y(N425) );
  INVX2TF U475 ( .A(N342), .Y(N338) );
  NOR2X1TF U476 ( .A(N101), .B(N342), .Y(N221) );
  NOR3X1TF U477 ( .A(N104), .B(N288), .C(N280), .Y(I_SCLK1) );
  NOR3X1TF U478 ( .A(\SCPU_CTRL_SPI_PUT_CNT_STATE[1] ), .B(N104), .C(N280), 
        .Y(I_SCLK2) );
  CLKBUFX2TF U479 ( .A(N296), .Y(N299) );
  INVX2TF U480 ( .A(I_CTRL_MODE[1]), .Y(N374) );
  OAI2BB1X1TF U481 ( .A0N(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[0] ), .A1N(
        \SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[1] ), .B0(N300), .Y(
        SCPU_CTRL_SPI_CCT_N51) );
  OAI2BB1X1TF U482 ( .A0N(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[2] ), .A1N(N300), 
        .B0(N301), .Y(SCPU_CTRL_SPI_CCT_N52) );
  OAI2BB1X1TF U483 ( .A0N(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[3] ), .A1N(N301), 
        .B0(N333), .Y(SCPU_CTRL_SPI_CCT_N53) );
  AO21X1TF U484 ( .A0(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[6] ), .A1(N302), .B0(
        N303), .Y(SCPU_CTRL_SPI_CCT_N56) );
  XOR2X1TF U485 ( .A(\SCPU_CTRL_SPI_CCT_CNT_BIT_LOAD[7] ), .B(N303), .Y(
        SCPU_CTRL_SPI_CCT_N57) );
  OAI221XLTF U486 ( .A0(N104), .A1(SCPU_CTRL_SPI_A_SPI[0]), .B0(N305), .B1(
        SCPU_CTRL_SPI_I_ADDR[0]), .C0(N327), .Y(N304) );
  NOR2BX1TF U487 ( .AN(SCPU_CTRL_SPI_CEN), .B(N327), .Y(CEN_AFTER_MUX) );
  AO22X1TF U488 ( .A0(N326), .A1(I_CTRL_SO), .B0(SCPU_CTRL_SPI_D_DATAOUT[0]), 
        .B1(N327), .Y(D_AFTER_MUX[0]) );
  AO22X1TF U489 ( .A0(N326), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[1] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[1]), .B1(N327), .Y(D_AFTER_MUX[1]) );
  AO22X1TF U490 ( .A0(N326), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[2] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[2]), .B1(N276), .Y(D_AFTER_MUX[2]) );
  AO22X1TF U491 ( .A0(N326), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[3] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[3]), .B1(N276), .Y(D_AFTER_MUX[3]) );
  AO22X1TF U492 ( .A0(N326), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[4] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[4]), .B1(N276), .Y(D_AFTER_MUX[4]) );
  AO22X1TF U493 ( .A0(N326), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[5] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[5]), .B1(N276), .Y(D_AFTER_MUX[5]) );
  AO22X1TF U494 ( .A0(N326), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[6] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[6]), .B1(N276), .Y(D_AFTER_MUX[6]) );
  AO22X1TF U495 ( .A0(N326), .A1(\SCPU_CTRL_SPI_CCT_REG_BITS[7] ), .B0(
        SCPU_CTRL_SPI_D_DATAOUT[7]), .B1(N276), .Y(D_AFTER_MUX[7]) );
  OAI221XLTF U496 ( .A0(N275), .A1(I_LOAD_N), .B0(N373), .B1(N329), .C0(
        I_CTRL_BGN), .Y(N328) );
  OAI2BB2XLTF U497 ( .B0(N373), .B1(N337), .A0N(N330), .A1N(N328), .Y(N216) );
  AO21X1TF U498 ( .A0(I_CTRL_MODE[0]), .A1(I_CTRL_MODE[1]), .B0(N335), .Y(N336) );
  NAND3X1TF U499 ( .A(N281), .B(N284), .C(N279), .Y(N430) );
  NAND3BX1TF U500 ( .AN(N430), .B(N282), .C(N285), .Y(N344) );
  OAI222X1TF U501 ( .A0(N429), .A1(N351), .B0(N346), .B1(N348), .C0(N283), 
        .C1(N345), .Y(N210) );
  NAND2X1TF U502 ( .A(N352), .B(N358), .Y(N354) );
  NAND3X1TF U503 ( .A(N361), .B(N355), .C(N354), .Y(N207) );
  NAND2X1TF U504 ( .A(N358), .B(N291), .Y(N357) );
  AO22X1TF U505 ( .A0(N371), .A1(SCPU_CTRL_SPI_PUT_SRAM_REGS[7]), .B0(
        Q_FROM_SRAM[7]), .B1(N370), .Y(N204) );
  AO22X1TF U506 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[0]), .B0(N271), .B1(I_ADC_PI[0]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[0]) );
  AO22X1TF U507 ( .A0(N272), .A1(SCPU_CTRL_SPI_FOUT[1]), .B0(N271), .B1(
        I_ADC_PI[1]), .Y(SCPU_CTRL_SPI_IO_DATAINA[1]) );
  AO22X1TF U508 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[2]), .B0(N271), .B1(I_ADC_PI[2]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[2]) );
  AO22X1TF U509 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[3]), .B0(N271), .B1(I_ADC_PI[3]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[3]) );
  AO22X1TF U510 ( .A0(\SCPU_CTRL_SPI_IO_CONTROL[5] ), .A1(
        SCPU_CTRL_SPI_FOUT[5]), .B0(N271), .B1(I_ADC_PI[5]), .Y(
        SCPU_CTRL_SPI_IO_DATAINA[5]) );
  OAI2BB2XLTF U511 ( .B0(N288), .B1(N280), .A0N(N288), .A1N(
        SCPU_CTRL_SPI_PUT_N106), .Y(SCPU_CTRL_SPI_PUT_N107) );
  NAND2X1TF U512 ( .A(N280), .B(N288), .Y(N396) );
  NAND3X1TF U513 ( .A(SCPU_CTRL_SPI_A_SPI[2]), .B(SCPU_CTRL_SPI_A_SPI[0]), .C(
        SCPU_CTRL_SPI_A_SPI[1]), .Y(N418) );
  NAND2X1TF U514 ( .A(N415), .B(SCPU_CTRL_SPI_A_SPI[3]), .Y(N414) );
  NOR2BX1TF U515 ( .AN(SCPU_CTRL_SPI_A_SPI[4]), .B(N414), .Y(N408) );
  NAND2X1TF U516 ( .A(N408), .B(SCPU_CTRL_SPI_A_SPI[5]), .Y(N407) );
  NOR2BX1TF U517 ( .AN(SCPU_CTRL_SPI_A_SPI[6]), .B(N407), .Y(N399) );
  NAND2BX1TF U518 ( .AN(N425), .B(N399), .Y(N402) );
  OAI2BB1X1TF U519 ( .A0N(N426), .A1N(N399), .B0(N273), .Y(N404) );
  AOI2BB2X1TF U520 ( .B0(\SCPU_CTRL_SPI_IO_DATAOUTA[7] ), .B1(N298), .A0N(
        SCPU_CTRL_SPI_A_SPI[7]), .A1N(N402), .Y(N403) );
endmodule

